//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.02
//Part Number: GW5AST-LV138FPG676AC2/I1
//Device: GW5AST-138B
//Device Version: B
//Created Time: Thu Apr 18 00:31:55 2024

module SRAM_SDPB (dout, clka, cea, clkb, ceb, oce, reset, ada, din, adb, byte_ena);

output [31:0] dout;
input clka;
input cea;
input clkb;
input ceb;
input oce;
input reset;
input [15:0] ada;
input [31:0] din;
input [15:0] adb;
input [3:0] byte_ena;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire lut_f_64;
wire lut_f_65;
wire lut_f_66;
wire lut_f_67;
wire lut_f_68;
wire lut_f_69;
wire lut_f_70;
wire lut_f_71;
wire lut_f_72;
wire lut_f_73;
wire lut_f_74;
wire lut_f_75;
wire lut_f_76;
wire lut_f_77;
wire lut_f_78;
wire lut_f_79;
wire lut_f_80;
wire lut_f_81;
wire lut_f_82;
wire lut_f_83;
wire lut_f_84;
wire lut_f_85;
wire lut_f_86;
wire lut_f_87;
wire lut_f_88;
wire lut_f_89;
wire lut_f_90;
wire lut_f_91;
wire lut_f_92;
wire lut_f_93;
wire lut_f_94;
wire lut_f_95;
wire lut_f_96;
wire lut_f_97;
wire lut_f_98;
wire lut_f_99;
wire lut_f_100;
wire lut_f_101;
wire lut_f_102;
wire lut_f_103;
wire lut_f_104;
wire lut_f_105;
wire lut_f_106;
wire lut_f_107;
wire lut_f_108;
wire lut_f_109;
wire lut_f_110;
wire lut_f_111;
wire lut_f_112;
wire lut_f_113;
wire lut_f_114;
wire lut_f_115;
wire lut_f_116;
wire lut_f_117;
wire lut_f_118;
wire lut_f_119;
wire lut_f_120;
wire lut_f_121;
wire lut_f_122;
wire lut_f_123;
wire lut_f_124;
wire lut_f_125;
wire lut_f_126;
wire lut_f_127;
wire [15:0] sdpb_inst_0_dout_w;
wire [15:0] sdpb_inst_0_dout;
wire [15:0] sdpb_inst_1_dout_w;
wire [15:0] sdpb_inst_1_dout;
wire [15:0] sdpb_inst_2_dout_w;
wire [15:0] sdpb_inst_2_dout;
wire [15:0] sdpb_inst_3_dout_w;
wire [15:0] sdpb_inst_3_dout;
wire [15:0] sdpb_inst_4_dout_w;
wire [15:0] sdpb_inst_4_dout;
wire [15:0] sdpb_inst_5_dout_w;
wire [15:0] sdpb_inst_5_dout;
wire [15:0] sdpb_inst_6_dout_w;
wire [15:0] sdpb_inst_6_dout;
wire [15:0] sdpb_inst_7_dout_w;
wire [15:0] sdpb_inst_7_dout;
wire [15:0] sdpb_inst_8_dout_w;
wire [15:0] sdpb_inst_8_dout;
wire [15:0] sdpb_inst_9_dout_w;
wire [15:0] sdpb_inst_9_dout;
wire [15:0] sdpb_inst_10_dout_w;
wire [15:0] sdpb_inst_10_dout;
wire [15:0] sdpb_inst_11_dout_w;
wire [15:0] sdpb_inst_11_dout;
wire [15:0] sdpb_inst_12_dout_w;
wire [15:0] sdpb_inst_12_dout;
wire [15:0] sdpb_inst_13_dout_w;
wire [15:0] sdpb_inst_13_dout;
wire [15:0] sdpb_inst_14_dout_w;
wire [15:0] sdpb_inst_14_dout;
wire [15:0] sdpb_inst_15_dout_w;
wire [15:0] sdpb_inst_15_dout;
wire [15:0] sdpb_inst_16_dout_w;
wire [15:0] sdpb_inst_16_dout;
wire [15:0] sdpb_inst_17_dout_w;
wire [15:0] sdpb_inst_17_dout;
wire [15:0] sdpb_inst_18_dout_w;
wire [15:0] sdpb_inst_18_dout;
wire [15:0] sdpb_inst_19_dout_w;
wire [15:0] sdpb_inst_19_dout;
wire [15:0] sdpb_inst_20_dout_w;
wire [15:0] sdpb_inst_20_dout;
wire [15:0] sdpb_inst_21_dout_w;
wire [15:0] sdpb_inst_21_dout;
wire [15:0] sdpb_inst_22_dout_w;
wire [15:0] sdpb_inst_22_dout;
wire [15:0] sdpb_inst_23_dout_w;
wire [15:0] sdpb_inst_23_dout;
wire [15:0] sdpb_inst_24_dout_w;
wire [15:0] sdpb_inst_24_dout;
wire [15:0] sdpb_inst_25_dout_w;
wire [15:0] sdpb_inst_25_dout;
wire [15:0] sdpb_inst_26_dout_w;
wire [15:0] sdpb_inst_26_dout;
wire [15:0] sdpb_inst_27_dout_w;
wire [15:0] sdpb_inst_27_dout;
wire [15:0] sdpb_inst_28_dout_w;
wire [15:0] sdpb_inst_28_dout;
wire [15:0] sdpb_inst_29_dout_w;
wire [15:0] sdpb_inst_29_dout;
wire [15:0] sdpb_inst_30_dout_w;
wire [15:0] sdpb_inst_30_dout;
wire [15:0] sdpb_inst_31_dout_w;
wire [15:0] sdpb_inst_31_dout;
wire [15:0] sdpb_inst_32_dout_w;
wire [15:0] sdpb_inst_32_dout;
wire [15:0] sdpb_inst_33_dout_w;
wire [15:0] sdpb_inst_33_dout;
wire [15:0] sdpb_inst_34_dout_w;
wire [15:0] sdpb_inst_34_dout;
wire [15:0] sdpb_inst_35_dout_w;
wire [15:0] sdpb_inst_35_dout;
wire [15:0] sdpb_inst_36_dout_w;
wire [15:0] sdpb_inst_36_dout;
wire [15:0] sdpb_inst_37_dout_w;
wire [15:0] sdpb_inst_37_dout;
wire [15:0] sdpb_inst_38_dout_w;
wire [15:0] sdpb_inst_38_dout;
wire [15:0] sdpb_inst_39_dout_w;
wire [15:0] sdpb_inst_39_dout;
wire [15:0] sdpb_inst_40_dout_w;
wire [15:0] sdpb_inst_40_dout;
wire [15:0] sdpb_inst_41_dout_w;
wire [15:0] sdpb_inst_41_dout;
wire [15:0] sdpb_inst_42_dout_w;
wire [15:0] sdpb_inst_42_dout;
wire [15:0] sdpb_inst_43_dout_w;
wire [15:0] sdpb_inst_43_dout;
wire [15:0] sdpb_inst_44_dout_w;
wire [15:0] sdpb_inst_44_dout;
wire [15:0] sdpb_inst_45_dout_w;
wire [15:0] sdpb_inst_45_dout;
wire [15:0] sdpb_inst_46_dout_w;
wire [15:0] sdpb_inst_46_dout;
wire [15:0] sdpb_inst_47_dout_w;
wire [15:0] sdpb_inst_47_dout;
wire [15:0] sdpb_inst_48_dout_w;
wire [15:0] sdpb_inst_48_dout;
wire [15:0] sdpb_inst_49_dout_w;
wire [15:0] sdpb_inst_49_dout;
wire [15:0] sdpb_inst_50_dout_w;
wire [15:0] sdpb_inst_50_dout;
wire [15:0] sdpb_inst_51_dout_w;
wire [15:0] sdpb_inst_51_dout;
wire [15:0] sdpb_inst_52_dout_w;
wire [15:0] sdpb_inst_52_dout;
wire [15:0] sdpb_inst_53_dout_w;
wire [15:0] sdpb_inst_53_dout;
wire [15:0] sdpb_inst_54_dout_w;
wire [15:0] sdpb_inst_54_dout;
wire [15:0] sdpb_inst_55_dout_w;
wire [15:0] sdpb_inst_55_dout;
wire [15:0] sdpb_inst_56_dout_w;
wire [15:0] sdpb_inst_56_dout;
wire [15:0] sdpb_inst_57_dout_w;
wire [15:0] sdpb_inst_57_dout;
wire [15:0] sdpb_inst_58_dout_w;
wire [15:0] sdpb_inst_58_dout;
wire [15:0] sdpb_inst_59_dout_w;
wire [15:0] sdpb_inst_59_dout;
wire [15:0] sdpb_inst_60_dout_w;
wire [15:0] sdpb_inst_60_dout;
wire [15:0] sdpb_inst_61_dout_w;
wire [15:0] sdpb_inst_61_dout;
wire [15:0] sdpb_inst_62_dout_w;
wire [15:0] sdpb_inst_62_dout;
wire [15:0] sdpb_inst_63_dout_w;
wire [15:0] sdpb_inst_63_dout;
wire [15:0] sdpb_inst_64_dout_w;
wire [31:16] sdpb_inst_64_dout;
wire [15:0] sdpb_inst_65_dout_w;
wire [31:16] sdpb_inst_65_dout;
wire [15:0] sdpb_inst_66_dout_w;
wire [31:16] sdpb_inst_66_dout;
wire [15:0] sdpb_inst_67_dout_w;
wire [31:16] sdpb_inst_67_dout;
wire [15:0] sdpb_inst_68_dout_w;
wire [31:16] sdpb_inst_68_dout;
wire [15:0] sdpb_inst_69_dout_w;
wire [31:16] sdpb_inst_69_dout;
wire [15:0] sdpb_inst_70_dout_w;
wire [31:16] sdpb_inst_70_dout;
wire [15:0] sdpb_inst_71_dout_w;
wire [31:16] sdpb_inst_71_dout;
wire [15:0] sdpb_inst_72_dout_w;
wire [31:16] sdpb_inst_72_dout;
wire [15:0] sdpb_inst_73_dout_w;
wire [31:16] sdpb_inst_73_dout;
wire [15:0] sdpb_inst_74_dout_w;
wire [31:16] sdpb_inst_74_dout;
wire [15:0] sdpb_inst_75_dout_w;
wire [31:16] sdpb_inst_75_dout;
wire [15:0] sdpb_inst_76_dout_w;
wire [31:16] sdpb_inst_76_dout;
wire [15:0] sdpb_inst_77_dout_w;
wire [31:16] sdpb_inst_77_dout;
wire [15:0] sdpb_inst_78_dout_w;
wire [31:16] sdpb_inst_78_dout;
wire [15:0] sdpb_inst_79_dout_w;
wire [31:16] sdpb_inst_79_dout;
wire [15:0] sdpb_inst_80_dout_w;
wire [31:16] sdpb_inst_80_dout;
wire [15:0] sdpb_inst_81_dout_w;
wire [31:16] sdpb_inst_81_dout;
wire [15:0] sdpb_inst_82_dout_w;
wire [31:16] sdpb_inst_82_dout;
wire [15:0] sdpb_inst_83_dout_w;
wire [31:16] sdpb_inst_83_dout;
wire [15:0] sdpb_inst_84_dout_w;
wire [31:16] sdpb_inst_84_dout;
wire [15:0] sdpb_inst_85_dout_w;
wire [31:16] sdpb_inst_85_dout;
wire [15:0] sdpb_inst_86_dout_w;
wire [31:16] sdpb_inst_86_dout;
wire [15:0] sdpb_inst_87_dout_w;
wire [31:16] sdpb_inst_87_dout;
wire [15:0] sdpb_inst_88_dout_w;
wire [31:16] sdpb_inst_88_dout;
wire [15:0] sdpb_inst_89_dout_w;
wire [31:16] sdpb_inst_89_dout;
wire [15:0] sdpb_inst_90_dout_w;
wire [31:16] sdpb_inst_90_dout;
wire [15:0] sdpb_inst_91_dout_w;
wire [31:16] sdpb_inst_91_dout;
wire [15:0] sdpb_inst_92_dout_w;
wire [31:16] sdpb_inst_92_dout;
wire [15:0] sdpb_inst_93_dout_w;
wire [31:16] sdpb_inst_93_dout;
wire [15:0] sdpb_inst_94_dout_w;
wire [31:16] sdpb_inst_94_dout;
wire [15:0] sdpb_inst_95_dout_w;
wire [31:16] sdpb_inst_95_dout;
wire [15:0] sdpb_inst_96_dout_w;
wire [31:16] sdpb_inst_96_dout;
wire [15:0] sdpb_inst_97_dout_w;
wire [31:16] sdpb_inst_97_dout;
wire [15:0] sdpb_inst_98_dout_w;
wire [31:16] sdpb_inst_98_dout;
wire [15:0] sdpb_inst_99_dout_w;
wire [31:16] sdpb_inst_99_dout;
wire [15:0] sdpb_inst_100_dout_w;
wire [31:16] sdpb_inst_100_dout;
wire [15:0] sdpb_inst_101_dout_w;
wire [31:16] sdpb_inst_101_dout;
wire [15:0] sdpb_inst_102_dout_w;
wire [31:16] sdpb_inst_102_dout;
wire [15:0] sdpb_inst_103_dout_w;
wire [31:16] sdpb_inst_103_dout;
wire [15:0] sdpb_inst_104_dout_w;
wire [31:16] sdpb_inst_104_dout;
wire [15:0] sdpb_inst_105_dout_w;
wire [31:16] sdpb_inst_105_dout;
wire [15:0] sdpb_inst_106_dout_w;
wire [31:16] sdpb_inst_106_dout;
wire [15:0] sdpb_inst_107_dout_w;
wire [31:16] sdpb_inst_107_dout;
wire [15:0] sdpb_inst_108_dout_w;
wire [31:16] sdpb_inst_108_dout;
wire [15:0] sdpb_inst_109_dout_w;
wire [31:16] sdpb_inst_109_dout;
wire [15:0] sdpb_inst_110_dout_w;
wire [31:16] sdpb_inst_110_dout;
wire [15:0] sdpb_inst_111_dout_w;
wire [31:16] sdpb_inst_111_dout;
wire [15:0] sdpb_inst_112_dout_w;
wire [31:16] sdpb_inst_112_dout;
wire [15:0] sdpb_inst_113_dout_w;
wire [31:16] sdpb_inst_113_dout;
wire [15:0] sdpb_inst_114_dout_w;
wire [31:16] sdpb_inst_114_dout;
wire [15:0] sdpb_inst_115_dout_w;
wire [31:16] sdpb_inst_115_dout;
wire [15:0] sdpb_inst_116_dout_w;
wire [31:16] sdpb_inst_116_dout;
wire [15:0] sdpb_inst_117_dout_w;
wire [31:16] sdpb_inst_117_dout;
wire [15:0] sdpb_inst_118_dout_w;
wire [31:16] sdpb_inst_118_dout;
wire [15:0] sdpb_inst_119_dout_w;
wire [31:16] sdpb_inst_119_dout;
wire [15:0] sdpb_inst_120_dout_w;
wire [31:16] sdpb_inst_120_dout;
wire [15:0] sdpb_inst_121_dout_w;
wire [31:16] sdpb_inst_121_dout;
wire [15:0] sdpb_inst_122_dout_w;
wire [31:16] sdpb_inst_122_dout;
wire [15:0] sdpb_inst_123_dout_w;
wire [31:16] sdpb_inst_123_dout;
wire [15:0] sdpb_inst_124_dout_w;
wire [31:16] sdpb_inst_124_dout;
wire [15:0] sdpb_inst_125_dout_w;
wire [31:16] sdpb_inst_125_dout;
wire [15:0] sdpb_inst_126_dout_w;
wire [31:16] sdpb_inst_126_dout;
wire [15:0] sdpb_inst_127_dout_w;
wire [31:16] sdpb_inst_127_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_588;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_867;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_888;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_898;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_929;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_960;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire mux_o_991;
wire mux_o_992;
wire mux_o_993;
wire mux_o_994;
wire mux_o_995;
wire mux_o_996;
wire mux_o_997;
wire mux_o_998;
wire mux_o_999;
wire mux_o_1000;
wire mux_o_1001;
wire mux_o_1002;
wire mux_o_1003;
wire mux_o_1004;
wire mux_o_1005;
wire mux_o_1006;
wire mux_o_1008;
wire mux_o_1009;
wire mux_o_1010;
wire mux_o_1011;
wire mux_o_1012;
wire mux_o_1013;
wire mux_o_1014;
wire mux_o_1015;
wire mux_o_1016;
wire mux_o_1017;
wire mux_o_1018;
wire mux_o_1019;
wire mux_o_1020;
wire mux_o_1021;
wire mux_o_1022;
wire mux_o_1023;
wire mux_o_1024;
wire mux_o_1025;
wire mux_o_1026;
wire mux_o_1027;
wire mux_o_1028;
wire mux_o_1029;
wire mux_o_1030;
wire mux_o_1031;
wire mux_o_1032;
wire mux_o_1033;
wire mux_o_1034;
wire mux_o_1035;
wire mux_o_1036;
wire mux_o_1037;
wire mux_o_1038;
wire mux_o_1039;
wire mux_o_1040;
wire mux_o_1041;
wire mux_o_1042;
wire mux_o_1043;
wire mux_o_1044;
wire mux_o_1045;
wire mux_o_1046;
wire mux_o_1047;
wire mux_o_1048;
wire mux_o_1049;
wire mux_o_1050;
wire mux_o_1051;
wire mux_o_1052;
wire mux_o_1053;
wire mux_o_1054;
wire mux_o_1055;
wire mux_o_1056;
wire mux_o_1057;
wire mux_o_1058;
wire mux_o_1059;
wire mux_o_1060;
wire mux_o_1061;
wire mux_o_1062;
wire mux_o_1063;
wire mux_o_1064;
wire mux_o_1065;
wire mux_o_1066;
wire mux_o_1067;
wire mux_o_1068;
wire mux_o_1069;
wire mux_o_1071;
wire mux_o_1072;
wire mux_o_1073;
wire mux_o_1074;
wire mux_o_1075;
wire mux_o_1076;
wire mux_o_1077;
wire mux_o_1078;
wire mux_o_1079;
wire mux_o_1080;
wire mux_o_1081;
wire mux_o_1082;
wire mux_o_1083;
wire mux_o_1084;
wire mux_o_1085;
wire mux_o_1086;
wire mux_o_1087;
wire mux_o_1088;
wire mux_o_1089;
wire mux_o_1090;
wire mux_o_1091;
wire mux_o_1092;
wire mux_o_1093;
wire mux_o_1094;
wire mux_o_1095;
wire mux_o_1096;
wire mux_o_1097;
wire mux_o_1098;
wire mux_o_1099;
wire mux_o_1100;
wire mux_o_1101;
wire mux_o_1102;
wire mux_o_1103;
wire mux_o_1104;
wire mux_o_1105;
wire mux_o_1106;
wire mux_o_1107;
wire mux_o_1108;
wire mux_o_1109;
wire mux_o_1110;
wire mux_o_1111;
wire mux_o_1112;
wire mux_o_1113;
wire mux_o_1114;
wire mux_o_1115;
wire mux_o_1116;
wire mux_o_1117;
wire mux_o_1118;
wire mux_o_1119;
wire mux_o_1120;
wire mux_o_1121;
wire mux_o_1122;
wire mux_o_1123;
wire mux_o_1124;
wire mux_o_1125;
wire mux_o_1126;
wire mux_o_1127;
wire mux_o_1128;
wire mux_o_1129;
wire mux_o_1130;
wire mux_o_1131;
wire mux_o_1132;
wire mux_o_1134;
wire mux_o_1135;
wire mux_o_1136;
wire mux_o_1137;
wire mux_o_1138;
wire mux_o_1139;
wire mux_o_1140;
wire mux_o_1141;
wire mux_o_1142;
wire mux_o_1143;
wire mux_o_1144;
wire mux_o_1145;
wire mux_o_1146;
wire mux_o_1147;
wire mux_o_1148;
wire mux_o_1149;
wire mux_o_1150;
wire mux_o_1151;
wire mux_o_1152;
wire mux_o_1153;
wire mux_o_1154;
wire mux_o_1155;
wire mux_o_1156;
wire mux_o_1157;
wire mux_o_1158;
wire mux_o_1159;
wire mux_o_1160;
wire mux_o_1161;
wire mux_o_1162;
wire mux_o_1163;
wire mux_o_1164;
wire mux_o_1165;
wire mux_o_1166;
wire mux_o_1167;
wire mux_o_1168;
wire mux_o_1169;
wire mux_o_1170;
wire mux_o_1171;
wire mux_o_1172;
wire mux_o_1173;
wire mux_o_1174;
wire mux_o_1175;
wire mux_o_1176;
wire mux_o_1177;
wire mux_o_1178;
wire mux_o_1179;
wire mux_o_1180;
wire mux_o_1181;
wire mux_o_1182;
wire mux_o_1183;
wire mux_o_1184;
wire mux_o_1185;
wire mux_o_1186;
wire mux_o_1187;
wire mux_o_1188;
wire mux_o_1189;
wire mux_o_1190;
wire mux_o_1191;
wire mux_o_1192;
wire mux_o_1193;
wire mux_o_1194;
wire mux_o_1195;
wire mux_o_1197;
wire mux_o_1198;
wire mux_o_1199;
wire mux_o_1200;
wire mux_o_1201;
wire mux_o_1202;
wire mux_o_1203;
wire mux_o_1204;
wire mux_o_1205;
wire mux_o_1206;
wire mux_o_1207;
wire mux_o_1208;
wire mux_o_1209;
wire mux_o_1210;
wire mux_o_1211;
wire mux_o_1212;
wire mux_o_1213;
wire mux_o_1214;
wire mux_o_1215;
wire mux_o_1216;
wire mux_o_1217;
wire mux_o_1218;
wire mux_o_1219;
wire mux_o_1220;
wire mux_o_1221;
wire mux_o_1222;
wire mux_o_1223;
wire mux_o_1224;
wire mux_o_1225;
wire mux_o_1226;
wire mux_o_1227;
wire mux_o_1228;
wire mux_o_1229;
wire mux_o_1230;
wire mux_o_1231;
wire mux_o_1232;
wire mux_o_1233;
wire mux_o_1234;
wire mux_o_1235;
wire mux_o_1236;
wire mux_o_1237;
wire mux_o_1238;
wire mux_o_1239;
wire mux_o_1240;
wire mux_o_1241;
wire mux_o_1242;
wire mux_o_1243;
wire mux_o_1244;
wire mux_o_1245;
wire mux_o_1246;
wire mux_o_1247;
wire mux_o_1248;
wire mux_o_1249;
wire mux_o_1250;
wire mux_o_1251;
wire mux_o_1252;
wire mux_o_1253;
wire mux_o_1254;
wire mux_o_1255;
wire mux_o_1256;
wire mux_o_1257;
wire mux_o_1258;
wire mux_o_1260;
wire mux_o_1261;
wire mux_o_1262;
wire mux_o_1263;
wire mux_o_1264;
wire mux_o_1265;
wire mux_o_1266;
wire mux_o_1267;
wire mux_o_1268;
wire mux_o_1269;
wire mux_o_1270;
wire mux_o_1271;
wire mux_o_1272;
wire mux_o_1273;
wire mux_o_1274;
wire mux_o_1275;
wire mux_o_1276;
wire mux_o_1277;
wire mux_o_1278;
wire mux_o_1279;
wire mux_o_1280;
wire mux_o_1281;
wire mux_o_1282;
wire mux_o_1283;
wire mux_o_1284;
wire mux_o_1285;
wire mux_o_1286;
wire mux_o_1287;
wire mux_o_1288;
wire mux_o_1289;
wire mux_o_1290;
wire mux_o_1291;
wire mux_o_1292;
wire mux_o_1293;
wire mux_o_1294;
wire mux_o_1295;
wire mux_o_1296;
wire mux_o_1297;
wire mux_o_1298;
wire mux_o_1299;
wire mux_o_1300;
wire mux_o_1301;
wire mux_o_1302;
wire mux_o_1303;
wire mux_o_1304;
wire mux_o_1305;
wire mux_o_1306;
wire mux_o_1307;
wire mux_o_1308;
wire mux_o_1309;
wire mux_o_1310;
wire mux_o_1311;
wire mux_o_1312;
wire mux_o_1313;
wire mux_o_1314;
wire mux_o_1315;
wire mux_o_1316;
wire mux_o_1317;
wire mux_o_1318;
wire mux_o_1319;
wire mux_o_1320;
wire mux_o_1321;
wire mux_o_1323;
wire mux_o_1324;
wire mux_o_1325;
wire mux_o_1326;
wire mux_o_1327;
wire mux_o_1328;
wire mux_o_1329;
wire mux_o_1330;
wire mux_o_1331;
wire mux_o_1332;
wire mux_o_1333;
wire mux_o_1334;
wire mux_o_1335;
wire mux_o_1336;
wire mux_o_1337;
wire mux_o_1338;
wire mux_o_1339;
wire mux_o_1340;
wire mux_o_1341;
wire mux_o_1342;
wire mux_o_1343;
wire mux_o_1344;
wire mux_o_1345;
wire mux_o_1346;
wire mux_o_1347;
wire mux_o_1348;
wire mux_o_1349;
wire mux_o_1350;
wire mux_o_1351;
wire mux_o_1352;
wire mux_o_1353;
wire mux_o_1354;
wire mux_o_1355;
wire mux_o_1356;
wire mux_o_1357;
wire mux_o_1358;
wire mux_o_1359;
wire mux_o_1360;
wire mux_o_1361;
wire mux_o_1362;
wire mux_o_1363;
wire mux_o_1364;
wire mux_o_1365;
wire mux_o_1366;
wire mux_o_1367;
wire mux_o_1368;
wire mux_o_1369;
wire mux_o_1370;
wire mux_o_1371;
wire mux_o_1372;
wire mux_o_1373;
wire mux_o_1374;
wire mux_o_1375;
wire mux_o_1376;
wire mux_o_1377;
wire mux_o_1378;
wire mux_o_1379;
wire mux_o_1380;
wire mux_o_1381;
wire mux_o_1382;
wire mux_o_1383;
wire mux_o_1384;
wire mux_o_1386;
wire mux_o_1387;
wire mux_o_1388;
wire mux_o_1389;
wire mux_o_1390;
wire mux_o_1391;
wire mux_o_1392;
wire mux_o_1393;
wire mux_o_1394;
wire mux_o_1395;
wire mux_o_1396;
wire mux_o_1397;
wire mux_o_1398;
wire mux_o_1399;
wire mux_o_1400;
wire mux_o_1401;
wire mux_o_1402;
wire mux_o_1403;
wire mux_o_1404;
wire mux_o_1405;
wire mux_o_1406;
wire mux_o_1407;
wire mux_o_1408;
wire mux_o_1409;
wire mux_o_1410;
wire mux_o_1411;
wire mux_o_1412;
wire mux_o_1413;
wire mux_o_1414;
wire mux_o_1415;
wire mux_o_1416;
wire mux_o_1417;
wire mux_o_1418;
wire mux_o_1419;
wire mux_o_1420;
wire mux_o_1421;
wire mux_o_1422;
wire mux_o_1423;
wire mux_o_1424;
wire mux_o_1425;
wire mux_o_1426;
wire mux_o_1427;
wire mux_o_1428;
wire mux_o_1429;
wire mux_o_1430;
wire mux_o_1431;
wire mux_o_1432;
wire mux_o_1433;
wire mux_o_1434;
wire mux_o_1435;
wire mux_o_1436;
wire mux_o_1437;
wire mux_o_1438;
wire mux_o_1439;
wire mux_o_1440;
wire mux_o_1441;
wire mux_o_1442;
wire mux_o_1443;
wire mux_o_1444;
wire mux_o_1445;
wire mux_o_1446;
wire mux_o_1447;
wire mux_o_1449;
wire mux_o_1450;
wire mux_o_1451;
wire mux_o_1452;
wire mux_o_1453;
wire mux_o_1454;
wire mux_o_1455;
wire mux_o_1456;
wire mux_o_1457;
wire mux_o_1458;
wire mux_o_1459;
wire mux_o_1460;
wire mux_o_1461;
wire mux_o_1462;
wire mux_o_1463;
wire mux_o_1464;
wire mux_o_1465;
wire mux_o_1466;
wire mux_o_1467;
wire mux_o_1468;
wire mux_o_1469;
wire mux_o_1470;
wire mux_o_1471;
wire mux_o_1472;
wire mux_o_1473;
wire mux_o_1474;
wire mux_o_1475;
wire mux_o_1476;
wire mux_o_1477;
wire mux_o_1478;
wire mux_o_1479;
wire mux_o_1480;
wire mux_o_1481;
wire mux_o_1482;
wire mux_o_1483;
wire mux_o_1484;
wire mux_o_1485;
wire mux_o_1486;
wire mux_o_1487;
wire mux_o_1488;
wire mux_o_1489;
wire mux_o_1490;
wire mux_o_1491;
wire mux_o_1492;
wire mux_o_1493;
wire mux_o_1494;
wire mux_o_1495;
wire mux_o_1496;
wire mux_o_1497;
wire mux_o_1498;
wire mux_o_1499;
wire mux_o_1500;
wire mux_o_1501;
wire mux_o_1502;
wire mux_o_1503;
wire mux_o_1504;
wire mux_o_1505;
wire mux_o_1506;
wire mux_o_1507;
wire mux_o_1508;
wire mux_o_1509;
wire mux_o_1510;
wire mux_o_1512;
wire mux_o_1513;
wire mux_o_1514;
wire mux_o_1515;
wire mux_o_1516;
wire mux_o_1517;
wire mux_o_1518;
wire mux_o_1519;
wire mux_o_1520;
wire mux_o_1521;
wire mux_o_1522;
wire mux_o_1523;
wire mux_o_1524;
wire mux_o_1525;
wire mux_o_1526;
wire mux_o_1527;
wire mux_o_1528;
wire mux_o_1529;
wire mux_o_1530;
wire mux_o_1531;
wire mux_o_1532;
wire mux_o_1533;
wire mux_o_1534;
wire mux_o_1535;
wire mux_o_1536;
wire mux_o_1537;
wire mux_o_1538;
wire mux_o_1539;
wire mux_o_1540;
wire mux_o_1541;
wire mux_o_1542;
wire mux_o_1543;
wire mux_o_1544;
wire mux_o_1545;
wire mux_o_1546;
wire mux_o_1547;
wire mux_o_1548;
wire mux_o_1549;
wire mux_o_1550;
wire mux_o_1551;
wire mux_o_1552;
wire mux_o_1553;
wire mux_o_1554;
wire mux_o_1555;
wire mux_o_1556;
wire mux_o_1557;
wire mux_o_1558;
wire mux_o_1559;
wire mux_o_1560;
wire mux_o_1561;
wire mux_o_1562;
wire mux_o_1563;
wire mux_o_1564;
wire mux_o_1565;
wire mux_o_1566;
wire mux_o_1567;
wire mux_o_1568;
wire mux_o_1569;
wire mux_o_1570;
wire mux_o_1571;
wire mux_o_1572;
wire mux_o_1573;
wire mux_o_1575;
wire mux_o_1576;
wire mux_o_1577;
wire mux_o_1578;
wire mux_o_1579;
wire mux_o_1580;
wire mux_o_1581;
wire mux_o_1582;
wire mux_o_1583;
wire mux_o_1584;
wire mux_o_1585;
wire mux_o_1586;
wire mux_o_1587;
wire mux_o_1588;
wire mux_o_1589;
wire mux_o_1590;
wire mux_o_1591;
wire mux_o_1592;
wire mux_o_1593;
wire mux_o_1594;
wire mux_o_1595;
wire mux_o_1596;
wire mux_o_1597;
wire mux_o_1598;
wire mux_o_1599;
wire mux_o_1600;
wire mux_o_1601;
wire mux_o_1602;
wire mux_o_1603;
wire mux_o_1604;
wire mux_o_1605;
wire mux_o_1606;
wire mux_o_1607;
wire mux_o_1608;
wire mux_o_1609;
wire mux_o_1610;
wire mux_o_1611;
wire mux_o_1612;
wire mux_o_1613;
wire mux_o_1614;
wire mux_o_1615;
wire mux_o_1616;
wire mux_o_1617;
wire mux_o_1618;
wire mux_o_1619;
wire mux_o_1620;
wire mux_o_1621;
wire mux_o_1622;
wire mux_o_1623;
wire mux_o_1624;
wire mux_o_1625;
wire mux_o_1626;
wire mux_o_1627;
wire mux_o_1628;
wire mux_o_1629;
wire mux_o_1630;
wire mux_o_1631;
wire mux_o_1632;
wire mux_o_1633;
wire mux_o_1634;
wire mux_o_1635;
wire mux_o_1636;
wire mux_o_1638;
wire mux_o_1639;
wire mux_o_1640;
wire mux_o_1641;
wire mux_o_1642;
wire mux_o_1643;
wire mux_o_1644;
wire mux_o_1645;
wire mux_o_1646;
wire mux_o_1647;
wire mux_o_1648;
wire mux_o_1649;
wire mux_o_1650;
wire mux_o_1651;
wire mux_o_1652;
wire mux_o_1653;
wire mux_o_1654;
wire mux_o_1655;
wire mux_o_1656;
wire mux_o_1657;
wire mux_o_1658;
wire mux_o_1659;
wire mux_o_1660;
wire mux_o_1661;
wire mux_o_1662;
wire mux_o_1663;
wire mux_o_1664;
wire mux_o_1665;
wire mux_o_1666;
wire mux_o_1667;
wire mux_o_1668;
wire mux_o_1669;
wire mux_o_1670;
wire mux_o_1671;
wire mux_o_1672;
wire mux_o_1673;
wire mux_o_1674;
wire mux_o_1675;
wire mux_o_1676;
wire mux_o_1677;
wire mux_o_1678;
wire mux_o_1679;
wire mux_o_1680;
wire mux_o_1681;
wire mux_o_1682;
wire mux_o_1683;
wire mux_o_1684;
wire mux_o_1685;
wire mux_o_1686;
wire mux_o_1687;
wire mux_o_1688;
wire mux_o_1689;
wire mux_o_1690;
wire mux_o_1691;
wire mux_o_1692;
wire mux_o_1693;
wire mux_o_1694;
wire mux_o_1695;
wire mux_o_1696;
wire mux_o_1697;
wire mux_o_1698;
wire mux_o_1699;
wire mux_o_1701;
wire mux_o_1702;
wire mux_o_1703;
wire mux_o_1704;
wire mux_o_1705;
wire mux_o_1706;
wire mux_o_1707;
wire mux_o_1708;
wire mux_o_1709;
wire mux_o_1710;
wire mux_o_1711;
wire mux_o_1712;
wire mux_o_1713;
wire mux_o_1714;
wire mux_o_1715;
wire mux_o_1716;
wire mux_o_1717;
wire mux_o_1718;
wire mux_o_1719;
wire mux_o_1720;
wire mux_o_1721;
wire mux_o_1722;
wire mux_o_1723;
wire mux_o_1724;
wire mux_o_1725;
wire mux_o_1726;
wire mux_o_1727;
wire mux_o_1728;
wire mux_o_1729;
wire mux_o_1730;
wire mux_o_1731;
wire mux_o_1732;
wire mux_o_1733;
wire mux_o_1734;
wire mux_o_1735;
wire mux_o_1736;
wire mux_o_1737;
wire mux_o_1738;
wire mux_o_1739;
wire mux_o_1740;
wire mux_o_1741;
wire mux_o_1742;
wire mux_o_1743;
wire mux_o_1744;
wire mux_o_1745;
wire mux_o_1746;
wire mux_o_1747;
wire mux_o_1748;
wire mux_o_1749;
wire mux_o_1750;
wire mux_o_1751;
wire mux_o_1752;
wire mux_o_1753;
wire mux_o_1754;
wire mux_o_1755;
wire mux_o_1756;
wire mux_o_1757;
wire mux_o_1758;
wire mux_o_1759;
wire mux_o_1760;
wire mux_o_1761;
wire mux_o_1762;
wire mux_o_1764;
wire mux_o_1765;
wire mux_o_1766;
wire mux_o_1767;
wire mux_o_1768;
wire mux_o_1769;
wire mux_o_1770;
wire mux_o_1771;
wire mux_o_1772;
wire mux_o_1773;
wire mux_o_1774;
wire mux_o_1775;
wire mux_o_1776;
wire mux_o_1777;
wire mux_o_1778;
wire mux_o_1779;
wire mux_o_1780;
wire mux_o_1781;
wire mux_o_1782;
wire mux_o_1783;
wire mux_o_1784;
wire mux_o_1785;
wire mux_o_1786;
wire mux_o_1787;
wire mux_o_1788;
wire mux_o_1789;
wire mux_o_1790;
wire mux_o_1791;
wire mux_o_1792;
wire mux_o_1793;
wire mux_o_1794;
wire mux_o_1795;
wire mux_o_1796;
wire mux_o_1797;
wire mux_o_1798;
wire mux_o_1799;
wire mux_o_1800;
wire mux_o_1801;
wire mux_o_1802;
wire mux_o_1803;
wire mux_o_1804;
wire mux_o_1805;
wire mux_o_1806;
wire mux_o_1807;
wire mux_o_1808;
wire mux_o_1809;
wire mux_o_1810;
wire mux_o_1811;
wire mux_o_1812;
wire mux_o_1813;
wire mux_o_1814;
wire mux_o_1815;
wire mux_o_1816;
wire mux_o_1817;
wire mux_o_1818;
wire mux_o_1819;
wire mux_o_1820;
wire mux_o_1821;
wire mux_o_1822;
wire mux_o_1823;
wire mux_o_1824;
wire mux_o_1825;
wire mux_o_1827;
wire mux_o_1828;
wire mux_o_1829;
wire mux_o_1830;
wire mux_o_1831;
wire mux_o_1832;
wire mux_o_1833;
wire mux_o_1834;
wire mux_o_1835;
wire mux_o_1836;
wire mux_o_1837;
wire mux_o_1838;
wire mux_o_1839;
wire mux_o_1840;
wire mux_o_1841;
wire mux_o_1842;
wire mux_o_1843;
wire mux_o_1844;
wire mux_o_1845;
wire mux_o_1846;
wire mux_o_1847;
wire mux_o_1848;
wire mux_o_1849;
wire mux_o_1850;
wire mux_o_1851;
wire mux_o_1852;
wire mux_o_1853;
wire mux_o_1854;
wire mux_o_1855;
wire mux_o_1856;
wire mux_o_1857;
wire mux_o_1858;
wire mux_o_1859;
wire mux_o_1860;
wire mux_o_1861;
wire mux_o_1862;
wire mux_o_1863;
wire mux_o_1864;
wire mux_o_1865;
wire mux_o_1866;
wire mux_o_1867;
wire mux_o_1868;
wire mux_o_1869;
wire mux_o_1870;
wire mux_o_1871;
wire mux_o_1872;
wire mux_o_1873;
wire mux_o_1874;
wire mux_o_1875;
wire mux_o_1876;
wire mux_o_1877;
wire mux_o_1878;
wire mux_o_1879;
wire mux_o_1880;
wire mux_o_1881;
wire mux_o_1882;
wire mux_o_1883;
wire mux_o_1884;
wire mux_o_1885;
wire mux_o_1886;
wire mux_o_1887;
wire mux_o_1888;
wire mux_o_1890;
wire mux_o_1891;
wire mux_o_1892;
wire mux_o_1893;
wire mux_o_1894;
wire mux_o_1895;
wire mux_o_1896;
wire mux_o_1897;
wire mux_o_1898;
wire mux_o_1899;
wire mux_o_1900;
wire mux_o_1901;
wire mux_o_1902;
wire mux_o_1903;
wire mux_o_1904;
wire mux_o_1905;
wire mux_o_1906;
wire mux_o_1907;
wire mux_o_1908;
wire mux_o_1909;
wire mux_o_1910;
wire mux_o_1911;
wire mux_o_1912;
wire mux_o_1913;
wire mux_o_1914;
wire mux_o_1915;
wire mux_o_1916;
wire mux_o_1917;
wire mux_o_1918;
wire mux_o_1919;
wire mux_o_1920;
wire mux_o_1921;
wire mux_o_1922;
wire mux_o_1923;
wire mux_o_1924;
wire mux_o_1925;
wire mux_o_1926;
wire mux_o_1927;
wire mux_o_1928;
wire mux_o_1929;
wire mux_o_1930;
wire mux_o_1931;
wire mux_o_1932;
wire mux_o_1933;
wire mux_o_1934;
wire mux_o_1935;
wire mux_o_1936;
wire mux_o_1937;
wire mux_o_1938;
wire mux_o_1939;
wire mux_o_1940;
wire mux_o_1941;
wire mux_o_1942;
wire mux_o_1943;
wire mux_o_1944;
wire mux_o_1945;
wire mux_o_1946;
wire mux_o_1947;
wire mux_o_1948;
wire mux_o_1949;
wire mux_o_1950;
wire mux_o_1951;
wire mux_o_1953;
wire mux_o_1954;
wire mux_o_1955;
wire mux_o_1956;
wire mux_o_1957;
wire mux_o_1958;
wire mux_o_1959;
wire mux_o_1960;
wire mux_o_1961;
wire mux_o_1962;
wire mux_o_1963;
wire mux_o_1964;
wire mux_o_1965;
wire mux_o_1966;
wire mux_o_1967;
wire mux_o_1968;
wire mux_o_1969;
wire mux_o_1970;
wire mux_o_1971;
wire mux_o_1972;
wire mux_o_1973;
wire mux_o_1974;
wire mux_o_1975;
wire mux_o_1976;
wire mux_o_1977;
wire mux_o_1978;
wire mux_o_1979;
wire mux_o_1980;
wire mux_o_1981;
wire mux_o_1982;
wire mux_o_1983;
wire mux_o_1984;
wire mux_o_1985;
wire mux_o_1986;
wire mux_o_1987;
wire mux_o_1988;
wire mux_o_1989;
wire mux_o_1990;
wire mux_o_1991;
wire mux_o_1992;
wire mux_o_1993;
wire mux_o_1994;
wire mux_o_1995;
wire mux_o_1996;
wire mux_o_1997;
wire mux_o_1998;
wire mux_o_1999;
wire mux_o_2000;
wire mux_o_2001;
wire mux_o_2002;
wire mux_o_2003;
wire mux_o_2004;
wire mux_o_2005;
wire mux_o_2006;
wire mux_o_2007;
wire mux_o_2008;
wire mux_o_2009;
wire mux_o_2010;
wire mux_o_2011;
wire mux_o_2012;
wire mux_o_2013;
wire mux_o_2014;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT6 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_0.INIT = 64'h0000000000000001;
LUT6 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_1.INIT = 64'h0000000000000002;
LUT6 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_2.INIT = 64'h0000000000000004;
LUT6 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_3.INIT = 64'h0000000000000008;
LUT6 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_4.INIT = 64'h0000000000000010;
LUT6 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_5.INIT = 64'h0000000000000020;
LUT6 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_6.INIT = 64'h0000000000000040;
LUT6 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_7.INIT = 64'h0000000000000080;
LUT6 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_8.INIT = 64'h0000000000000100;
LUT6 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_9.INIT = 64'h0000000000000200;
LUT6 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_10.INIT = 64'h0000000000000400;
LUT6 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_11.INIT = 64'h0000000000000800;
LUT6 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_12.INIT = 64'h0000000000001000;
LUT6 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_13.INIT = 64'h0000000000002000;
LUT6 lut_inst_14 (
  .F(lut_f_14),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_14.INIT = 64'h0000000000004000;
LUT6 lut_inst_15 (
  .F(lut_f_15),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_15.INIT = 64'h0000000000008000;
LUT6 lut_inst_16 (
  .F(lut_f_16),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_16.INIT = 64'h0000000000010000;
LUT6 lut_inst_17 (
  .F(lut_f_17),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_17.INIT = 64'h0000000000020000;
LUT6 lut_inst_18 (
  .F(lut_f_18),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_18.INIT = 64'h0000000000040000;
LUT6 lut_inst_19 (
  .F(lut_f_19),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_19.INIT = 64'h0000000000080000;
LUT6 lut_inst_20 (
  .F(lut_f_20),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_20.INIT = 64'h0000000000100000;
LUT6 lut_inst_21 (
  .F(lut_f_21),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_21.INIT = 64'h0000000000200000;
LUT6 lut_inst_22 (
  .F(lut_f_22),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_22.INIT = 64'h0000000000400000;
LUT6 lut_inst_23 (
  .F(lut_f_23),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_23.INIT = 64'h0000000000800000;
LUT6 lut_inst_24 (
  .F(lut_f_24),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_24.INIT = 64'h0000000001000000;
LUT6 lut_inst_25 (
  .F(lut_f_25),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_25.INIT = 64'h0000000002000000;
LUT6 lut_inst_26 (
  .F(lut_f_26),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_26.INIT = 64'h0000000004000000;
LUT6 lut_inst_27 (
  .F(lut_f_27),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_27.INIT = 64'h0000000008000000;
LUT6 lut_inst_28 (
  .F(lut_f_28),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_28.INIT = 64'h0000000010000000;
LUT6 lut_inst_29 (
  .F(lut_f_29),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_29.INIT = 64'h0000000020000000;
LUT6 lut_inst_30 (
  .F(lut_f_30),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_30.INIT = 64'h0000000040000000;
LUT6 lut_inst_31 (
  .F(lut_f_31),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_31.INIT = 64'h0000000080000000;
LUT6 lut_inst_32 (
  .F(lut_f_32),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_32.INIT = 64'h0000000100000000;
LUT6 lut_inst_33 (
  .F(lut_f_33),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_33.INIT = 64'h0000000200000000;
LUT6 lut_inst_34 (
  .F(lut_f_34),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_34.INIT = 64'h0000000400000000;
LUT6 lut_inst_35 (
  .F(lut_f_35),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_35.INIT = 64'h0000000800000000;
LUT6 lut_inst_36 (
  .F(lut_f_36),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_36.INIT = 64'h0000001000000000;
LUT6 lut_inst_37 (
  .F(lut_f_37),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_37.INIT = 64'h0000002000000000;
LUT6 lut_inst_38 (
  .F(lut_f_38),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_38.INIT = 64'h0000004000000000;
LUT6 lut_inst_39 (
  .F(lut_f_39),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_39.INIT = 64'h0000008000000000;
LUT6 lut_inst_40 (
  .F(lut_f_40),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_40.INIT = 64'h0000010000000000;
LUT6 lut_inst_41 (
  .F(lut_f_41),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_41.INIT = 64'h0000020000000000;
LUT6 lut_inst_42 (
  .F(lut_f_42),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_42.INIT = 64'h0000040000000000;
LUT6 lut_inst_43 (
  .F(lut_f_43),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_43.INIT = 64'h0000080000000000;
LUT6 lut_inst_44 (
  .F(lut_f_44),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_44.INIT = 64'h0000100000000000;
LUT6 lut_inst_45 (
  .F(lut_f_45),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_45.INIT = 64'h0000200000000000;
LUT6 lut_inst_46 (
  .F(lut_f_46),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_46.INIT = 64'h0000400000000000;
LUT6 lut_inst_47 (
  .F(lut_f_47),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_47.INIT = 64'h0000800000000000;
LUT6 lut_inst_48 (
  .F(lut_f_48),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_48.INIT = 64'h0001000000000000;
LUT6 lut_inst_49 (
  .F(lut_f_49),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_49.INIT = 64'h0002000000000000;
LUT6 lut_inst_50 (
  .F(lut_f_50),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_50.INIT = 64'h0004000000000000;
LUT6 lut_inst_51 (
  .F(lut_f_51),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_51.INIT = 64'h0008000000000000;
LUT6 lut_inst_52 (
  .F(lut_f_52),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_52.INIT = 64'h0010000000000000;
LUT6 lut_inst_53 (
  .F(lut_f_53),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_53.INIT = 64'h0020000000000000;
LUT6 lut_inst_54 (
  .F(lut_f_54),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_54.INIT = 64'h0040000000000000;
LUT6 lut_inst_55 (
  .F(lut_f_55),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_55.INIT = 64'h0080000000000000;
LUT6 lut_inst_56 (
  .F(lut_f_56),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_56.INIT = 64'h0100000000000000;
LUT6 lut_inst_57 (
  .F(lut_f_57),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_57.INIT = 64'h0200000000000000;
LUT6 lut_inst_58 (
  .F(lut_f_58),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_58.INIT = 64'h0400000000000000;
LUT6 lut_inst_59 (
  .F(lut_f_59),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_59.INIT = 64'h0800000000000000;
LUT6 lut_inst_60 (
  .F(lut_f_60),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_60.INIT = 64'h1000000000000000;
LUT6 lut_inst_61 (
  .F(lut_f_61),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_61.INIT = 64'h2000000000000000;
LUT6 lut_inst_62 (
  .F(lut_f_62),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_62.INIT = 64'h4000000000000000;
LUT6 lut_inst_63 (
  .F(lut_f_63),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15])
);
defparam lut_inst_63.INIT = 64'h8000000000000000;
LUT6 lut_inst_64 (
  .F(lut_f_64),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_64.INIT = 64'h0000000000000001;
LUT6 lut_inst_65 (
  .F(lut_f_65),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_65.INIT = 64'h0000000000000002;
LUT6 lut_inst_66 (
  .F(lut_f_66),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_66.INIT = 64'h0000000000000004;
LUT6 lut_inst_67 (
  .F(lut_f_67),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_67.INIT = 64'h0000000000000008;
LUT6 lut_inst_68 (
  .F(lut_f_68),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_68.INIT = 64'h0000000000000010;
LUT6 lut_inst_69 (
  .F(lut_f_69),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_69.INIT = 64'h0000000000000020;
LUT6 lut_inst_70 (
  .F(lut_f_70),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_70.INIT = 64'h0000000000000040;
LUT6 lut_inst_71 (
  .F(lut_f_71),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_71.INIT = 64'h0000000000000080;
LUT6 lut_inst_72 (
  .F(lut_f_72),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_72.INIT = 64'h0000000000000100;
LUT6 lut_inst_73 (
  .F(lut_f_73),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_73.INIT = 64'h0000000000000200;
LUT6 lut_inst_74 (
  .F(lut_f_74),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_74.INIT = 64'h0000000000000400;
LUT6 lut_inst_75 (
  .F(lut_f_75),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_75.INIT = 64'h0000000000000800;
LUT6 lut_inst_76 (
  .F(lut_f_76),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_76.INIT = 64'h0000000000001000;
LUT6 lut_inst_77 (
  .F(lut_f_77),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_77.INIT = 64'h0000000000002000;
LUT6 lut_inst_78 (
  .F(lut_f_78),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_78.INIT = 64'h0000000000004000;
LUT6 lut_inst_79 (
  .F(lut_f_79),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_79.INIT = 64'h0000000000008000;
LUT6 lut_inst_80 (
  .F(lut_f_80),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_80.INIT = 64'h0000000000010000;
LUT6 lut_inst_81 (
  .F(lut_f_81),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_81.INIT = 64'h0000000000020000;
LUT6 lut_inst_82 (
  .F(lut_f_82),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_82.INIT = 64'h0000000000040000;
LUT6 lut_inst_83 (
  .F(lut_f_83),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_83.INIT = 64'h0000000000080000;
LUT6 lut_inst_84 (
  .F(lut_f_84),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_84.INIT = 64'h0000000000100000;
LUT6 lut_inst_85 (
  .F(lut_f_85),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_85.INIT = 64'h0000000000200000;
LUT6 lut_inst_86 (
  .F(lut_f_86),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_86.INIT = 64'h0000000000400000;
LUT6 lut_inst_87 (
  .F(lut_f_87),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_87.INIT = 64'h0000000000800000;
LUT6 lut_inst_88 (
  .F(lut_f_88),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_88.INIT = 64'h0000000001000000;
LUT6 lut_inst_89 (
  .F(lut_f_89),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_89.INIT = 64'h0000000002000000;
LUT6 lut_inst_90 (
  .F(lut_f_90),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_90.INIT = 64'h0000000004000000;
LUT6 lut_inst_91 (
  .F(lut_f_91),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_91.INIT = 64'h0000000008000000;
LUT6 lut_inst_92 (
  .F(lut_f_92),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_92.INIT = 64'h0000000010000000;
LUT6 lut_inst_93 (
  .F(lut_f_93),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_93.INIT = 64'h0000000020000000;
LUT6 lut_inst_94 (
  .F(lut_f_94),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_94.INIT = 64'h0000000040000000;
LUT6 lut_inst_95 (
  .F(lut_f_95),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_95.INIT = 64'h0000000080000000;
LUT6 lut_inst_96 (
  .F(lut_f_96),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_96.INIT = 64'h0000000100000000;
LUT6 lut_inst_97 (
  .F(lut_f_97),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_97.INIT = 64'h0000000200000000;
LUT6 lut_inst_98 (
  .F(lut_f_98),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_98.INIT = 64'h0000000400000000;
LUT6 lut_inst_99 (
  .F(lut_f_99),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_99.INIT = 64'h0000000800000000;
LUT6 lut_inst_100 (
  .F(lut_f_100),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_100.INIT = 64'h0000001000000000;
LUT6 lut_inst_101 (
  .F(lut_f_101),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_101.INIT = 64'h0000002000000000;
LUT6 lut_inst_102 (
  .F(lut_f_102),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_102.INIT = 64'h0000004000000000;
LUT6 lut_inst_103 (
  .F(lut_f_103),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_103.INIT = 64'h0000008000000000;
LUT6 lut_inst_104 (
  .F(lut_f_104),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_104.INIT = 64'h0000010000000000;
LUT6 lut_inst_105 (
  .F(lut_f_105),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_105.INIT = 64'h0000020000000000;
LUT6 lut_inst_106 (
  .F(lut_f_106),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_106.INIT = 64'h0000040000000000;
LUT6 lut_inst_107 (
  .F(lut_f_107),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_107.INIT = 64'h0000080000000000;
LUT6 lut_inst_108 (
  .F(lut_f_108),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_108.INIT = 64'h0000100000000000;
LUT6 lut_inst_109 (
  .F(lut_f_109),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_109.INIT = 64'h0000200000000000;
LUT6 lut_inst_110 (
  .F(lut_f_110),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_110.INIT = 64'h0000400000000000;
LUT6 lut_inst_111 (
  .F(lut_f_111),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_111.INIT = 64'h0000800000000000;
LUT6 lut_inst_112 (
  .F(lut_f_112),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_112.INIT = 64'h0001000000000000;
LUT6 lut_inst_113 (
  .F(lut_f_113),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_113.INIT = 64'h0002000000000000;
LUT6 lut_inst_114 (
  .F(lut_f_114),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_114.INIT = 64'h0004000000000000;
LUT6 lut_inst_115 (
  .F(lut_f_115),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_115.INIT = 64'h0008000000000000;
LUT6 lut_inst_116 (
  .F(lut_f_116),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_116.INIT = 64'h0010000000000000;
LUT6 lut_inst_117 (
  .F(lut_f_117),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_117.INIT = 64'h0020000000000000;
LUT6 lut_inst_118 (
  .F(lut_f_118),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_118.INIT = 64'h0040000000000000;
LUT6 lut_inst_119 (
  .F(lut_f_119),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_119.INIT = 64'h0080000000000000;
LUT6 lut_inst_120 (
  .F(lut_f_120),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_120.INIT = 64'h0100000000000000;
LUT6 lut_inst_121 (
  .F(lut_f_121),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_121.INIT = 64'h0200000000000000;
LUT6 lut_inst_122 (
  .F(lut_f_122),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_122.INIT = 64'h0400000000000000;
LUT6 lut_inst_123 (
  .F(lut_f_123),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_123.INIT = 64'h0800000000000000;
LUT6 lut_inst_124 (
  .F(lut_f_124),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_124.INIT = 64'h1000000000000000;
LUT6 lut_inst_125 (
  .F(lut_f_125),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_125.INIT = 64'h2000000000000000;
LUT6 lut_inst_126 (
  .F(lut_f_126),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_126.INIT = 64'h4000000000000000;
LUT6 lut_inst_127 (
  .F(lut_f_127),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15])
);
defparam lut_inst_127.INIT = 64'h8000000000000000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],sdpb_inst_0_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_64}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_0.RESET_MODE = "SYNC";

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[15:0],sdpb_inst_1_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_65}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 16;
defparam sdpb_inst_1.BIT_WIDTH_1 = 16;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[15:0],sdpb_inst_2_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_66}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 16;
defparam sdpb_inst_2.BIT_WIDTH_1 = 16;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_2.RESET_MODE = "SYNC";

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[15:0],sdpb_inst_3_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_67}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 16;
defparam sdpb_inst_3.BIT_WIDTH_1 = 16;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[15:0],sdpb_inst_4_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_68}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 16;
defparam sdpb_inst_4.BIT_WIDTH_1 = 16;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_4.RESET_MODE = "SYNC";

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[15:0],sdpb_inst_5_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_69}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 16;
defparam sdpb_inst_5.BIT_WIDTH_1 = 16;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[15:0],sdpb_inst_6_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_70}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 16;
defparam sdpb_inst_6.BIT_WIDTH_1 = 16;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_6.RESET_MODE = "SYNC";

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[15:0],sdpb_inst_7_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_71}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 16;
defparam sdpb_inst_7.BIT_WIDTH_1 = 16;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[15:0],sdpb_inst_8_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_72}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 16;
defparam sdpb_inst_8.BIT_WIDTH_1 = 16;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[15:0],sdpb_inst_9_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_73}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_9.READ_MODE = 1'b0;
defparam sdpb_inst_9.BIT_WIDTH_0 = 16;
defparam sdpb_inst_9.BIT_WIDTH_1 = 16;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_9.RESET_MODE = "SYNC";

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[15:0],sdpb_inst_10_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_74}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_10.READ_MODE = 1'b0;
defparam sdpb_inst_10.BIT_WIDTH_0 = 16;
defparam sdpb_inst_10.BIT_WIDTH_1 = 16;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_10.RESET_MODE = "SYNC";

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[15:0],sdpb_inst_11_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_75}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_11.READ_MODE = 1'b0;
defparam sdpb_inst_11.BIT_WIDTH_0 = 16;
defparam sdpb_inst_11.BIT_WIDTH_1 = 16;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_11.RESET_MODE = "SYNC";

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[15:0],sdpb_inst_12_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_76}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_12.READ_MODE = 1'b0;
defparam sdpb_inst_12.BIT_WIDTH_0 = 16;
defparam sdpb_inst_12.BIT_WIDTH_1 = 16;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_12.RESET_MODE = "SYNC";

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[15:0],sdpb_inst_13_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_77}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_13.READ_MODE = 1'b0;
defparam sdpb_inst_13.BIT_WIDTH_0 = 16;
defparam sdpb_inst_13.BIT_WIDTH_1 = 16;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_13.RESET_MODE = "SYNC";

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[15:0],sdpb_inst_14_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_78}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_14.READ_MODE = 1'b0;
defparam sdpb_inst_14.BIT_WIDTH_0 = 16;
defparam sdpb_inst_14.BIT_WIDTH_1 = 16;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_14.RESET_MODE = "SYNC";

SDPB sdpb_inst_15 (
    .DO({sdpb_inst_15_dout_w[15:0],sdpb_inst_15_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_79}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_15.READ_MODE = 1'b0;
defparam sdpb_inst_15.BIT_WIDTH_0 = 16;
defparam sdpb_inst_15.BIT_WIDTH_1 = 16;
defparam sdpb_inst_15.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_15.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_15.RESET_MODE = "SYNC";

SDPB sdpb_inst_16 (
    .DO({sdpb_inst_16_dout_w[15:0],sdpb_inst_16_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_16}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_80}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_16.READ_MODE = 1'b0;
defparam sdpb_inst_16.BIT_WIDTH_0 = 16;
defparam sdpb_inst_16.BIT_WIDTH_1 = 16;
defparam sdpb_inst_16.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_16.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_16.RESET_MODE = "SYNC";

SDPB sdpb_inst_17 (
    .DO({sdpb_inst_17_dout_w[15:0],sdpb_inst_17_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_17}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_81}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_17.READ_MODE = 1'b0;
defparam sdpb_inst_17.BIT_WIDTH_0 = 16;
defparam sdpb_inst_17.BIT_WIDTH_1 = 16;
defparam sdpb_inst_17.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_17.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_17.RESET_MODE = "SYNC";

SDPB sdpb_inst_18 (
    .DO({sdpb_inst_18_dout_w[15:0],sdpb_inst_18_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_18}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_82}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_18.READ_MODE = 1'b0;
defparam sdpb_inst_18.BIT_WIDTH_0 = 16;
defparam sdpb_inst_18.BIT_WIDTH_1 = 16;
defparam sdpb_inst_18.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_18.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_18.RESET_MODE = "SYNC";

SDPB sdpb_inst_19 (
    .DO({sdpb_inst_19_dout_w[15:0],sdpb_inst_19_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_19}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_83}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_19.READ_MODE = 1'b0;
defparam sdpb_inst_19.BIT_WIDTH_0 = 16;
defparam sdpb_inst_19.BIT_WIDTH_1 = 16;
defparam sdpb_inst_19.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_19.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_19.RESET_MODE = "SYNC";

SDPB sdpb_inst_20 (
    .DO({sdpb_inst_20_dout_w[15:0],sdpb_inst_20_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_20}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_84}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_20.READ_MODE = 1'b0;
defparam sdpb_inst_20.BIT_WIDTH_0 = 16;
defparam sdpb_inst_20.BIT_WIDTH_1 = 16;
defparam sdpb_inst_20.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_20.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_20.RESET_MODE = "SYNC";

SDPB sdpb_inst_21 (
    .DO({sdpb_inst_21_dout_w[15:0],sdpb_inst_21_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_21}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_85}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_21.READ_MODE = 1'b0;
defparam sdpb_inst_21.BIT_WIDTH_0 = 16;
defparam sdpb_inst_21.BIT_WIDTH_1 = 16;
defparam sdpb_inst_21.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_21.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_21.RESET_MODE = "SYNC";

SDPB sdpb_inst_22 (
    .DO({sdpb_inst_22_dout_w[15:0],sdpb_inst_22_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_22}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_86}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_22.READ_MODE = 1'b0;
defparam sdpb_inst_22.BIT_WIDTH_0 = 16;
defparam sdpb_inst_22.BIT_WIDTH_1 = 16;
defparam sdpb_inst_22.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_22.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_22.RESET_MODE = "SYNC";

SDPB sdpb_inst_23 (
    .DO({sdpb_inst_23_dout_w[15:0],sdpb_inst_23_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_23}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_87}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_23.READ_MODE = 1'b0;
defparam sdpb_inst_23.BIT_WIDTH_0 = 16;
defparam sdpb_inst_23.BIT_WIDTH_1 = 16;
defparam sdpb_inst_23.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_23.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_23.RESET_MODE = "SYNC";

SDPB sdpb_inst_24 (
    .DO({sdpb_inst_24_dout_w[15:0],sdpb_inst_24_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_24}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_88}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_24.READ_MODE = 1'b0;
defparam sdpb_inst_24.BIT_WIDTH_0 = 16;
defparam sdpb_inst_24.BIT_WIDTH_1 = 16;
defparam sdpb_inst_24.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_24.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_24.RESET_MODE = "SYNC";

SDPB sdpb_inst_25 (
    .DO({sdpb_inst_25_dout_w[15:0],sdpb_inst_25_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_25}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_89}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_25.READ_MODE = 1'b0;
defparam sdpb_inst_25.BIT_WIDTH_0 = 16;
defparam sdpb_inst_25.BIT_WIDTH_1 = 16;
defparam sdpb_inst_25.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_25.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_25.RESET_MODE = "SYNC";

SDPB sdpb_inst_26 (
    .DO({sdpb_inst_26_dout_w[15:0],sdpb_inst_26_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_26}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_90}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_26.READ_MODE = 1'b0;
defparam sdpb_inst_26.BIT_WIDTH_0 = 16;
defparam sdpb_inst_26.BIT_WIDTH_1 = 16;
defparam sdpb_inst_26.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_26.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_26.RESET_MODE = "SYNC";

SDPB sdpb_inst_27 (
    .DO({sdpb_inst_27_dout_w[15:0],sdpb_inst_27_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_27}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_91}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_27.READ_MODE = 1'b0;
defparam sdpb_inst_27.BIT_WIDTH_0 = 16;
defparam sdpb_inst_27.BIT_WIDTH_1 = 16;
defparam sdpb_inst_27.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_27.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_27.RESET_MODE = "SYNC";

SDPB sdpb_inst_28 (
    .DO({sdpb_inst_28_dout_w[15:0],sdpb_inst_28_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_28}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_92}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_28.READ_MODE = 1'b0;
defparam sdpb_inst_28.BIT_WIDTH_0 = 16;
defparam sdpb_inst_28.BIT_WIDTH_1 = 16;
defparam sdpb_inst_28.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_28.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_28.RESET_MODE = "SYNC";

SDPB sdpb_inst_29 (
    .DO({sdpb_inst_29_dout_w[15:0],sdpb_inst_29_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_29}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_93}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_29.READ_MODE = 1'b0;
defparam sdpb_inst_29.BIT_WIDTH_0 = 16;
defparam sdpb_inst_29.BIT_WIDTH_1 = 16;
defparam sdpb_inst_29.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_29.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_29.RESET_MODE = "SYNC";

SDPB sdpb_inst_30 (
    .DO({sdpb_inst_30_dout_w[15:0],sdpb_inst_30_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_30}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_94}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_30.READ_MODE = 1'b0;
defparam sdpb_inst_30.BIT_WIDTH_0 = 16;
defparam sdpb_inst_30.BIT_WIDTH_1 = 16;
defparam sdpb_inst_30.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_30.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_30.RESET_MODE = "SYNC";

SDPB sdpb_inst_31 (
    .DO({sdpb_inst_31_dout_w[15:0],sdpb_inst_31_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_31}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_95}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_31.READ_MODE = 1'b0;
defparam sdpb_inst_31.BIT_WIDTH_0 = 16;
defparam sdpb_inst_31.BIT_WIDTH_1 = 16;
defparam sdpb_inst_31.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_31.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_31.RESET_MODE = "SYNC";

SDPB sdpb_inst_32 (
    .DO({sdpb_inst_32_dout_w[15:0],sdpb_inst_32_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_32}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_96}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_32.READ_MODE = 1'b0;
defparam sdpb_inst_32.BIT_WIDTH_0 = 16;
defparam sdpb_inst_32.BIT_WIDTH_1 = 16;
defparam sdpb_inst_32.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_32.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_32.RESET_MODE = "SYNC";

SDPB sdpb_inst_33 (
    .DO({sdpb_inst_33_dout_w[15:0],sdpb_inst_33_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_33}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_97}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_33.READ_MODE = 1'b0;
defparam sdpb_inst_33.BIT_WIDTH_0 = 16;
defparam sdpb_inst_33.BIT_WIDTH_1 = 16;
defparam sdpb_inst_33.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_33.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_33.RESET_MODE = "SYNC";

SDPB sdpb_inst_34 (
    .DO({sdpb_inst_34_dout_w[15:0],sdpb_inst_34_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_34}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_98}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_34.READ_MODE = 1'b0;
defparam sdpb_inst_34.BIT_WIDTH_0 = 16;
defparam sdpb_inst_34.BIT_WIDTH_1 = 16;
defparam sdpb_inst_34.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_34.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_34.RESET_MODE = "SYNC";

SDPB sdpb_inst_35 (
    .DO({sdpb_inst_35_dout_w[15:0],sdpb_inst_35_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_35}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_99}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_35.READ_MODE = 1'b0;
defparam sdpb_inst_35.BIT_WIDTH_0 = 16;
defparam sdpb_inst_35.BIT_WIDTH_1 = 16;
defparam sdpb_inst_35.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_35.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_35.RESET_MODE = "SYNC";

SDPB sdpb_inst_36 (
    .DO({sdpb_inst_36_dout_w[15:0],sdpb_inst_36_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_36}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_100}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_36.READ_MODE = 1'b0;
defparam sdpb_inst_36.BIT_WIDTH_0 = 16;
defparam sdpb_inst_36.BIT_WIDTH_1 = 16;
defparam sdpb_inst_36.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_36.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_36.RESET_MODE = "SYNC";

SDPB sdpb_inst_37 (
    .DO({sdpb_inst_37_dout_w[15:0],sdpb_inst_37_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_37}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_101}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_37.READ_MODE = 1'b0;
defparam sdpb_inst_37.BIT_WIDTH_0 = 16;
defparam sdpb_inst_37.BIT_WIDTH_1 = 16;
defparam sdpb_inst_37.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_37.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_37.RESET_MODE = "SYNC";

SDPB sdpb_inst_38 (
    .DO({sdpb_inst_38_dout_w[15:0],sdpb_inst_38_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_38}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_102}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_38.READ_MODE = 1'b0;
defparam sdpb_inst_38.BIT_WIDTH_0 = 16;
defparam sdpb_inst_38.BIT_WIDTH_1 = 16;
defparam sdpb_inst_38.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_38.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_38.RESET_MODE = "SYNC";

SDPB sdpb_inst_39 (
    .DO({sdpb_inst_39_dout_w[15:0],sdpb_inst_39_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_39}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_103}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_39.READ_MODE = 1'b0;
defparam sdpb_inst_39.BIT_WIDTH_0 = 16;
defparam sdpb_inst_39.BIT_WIDTH_1 = 16;
defparam sdpb_inst_39.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_39.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_39.RESET_MODE = "SYNC";

SDPB sdpb_inst_40 (
    .DO({sdpb_inst_40_dout_w[15:0],sdpb_inst_40_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_40}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_104}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_40.READ_MODE = 1'b0;
defparam sdpb_inst_40.BIT_WIDTH_0 = 16;
defparam sdpb_inst_40.BIT_WIDTH_1 = 16;
defparam sdpb_inst_40.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_40.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_40.RESET_MODE = "SYNC";

SDPB sdpb_inst_41 (
    .DO({sdpb_inst_41_dout_w[15:0],sdpb_inst_41_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_41}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_105}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_41.READ_MODE = 1'b0;
defparam sdpb_inst_41.BIT_WIDTH_0 = 16;
defparam sdpb_inst_41.BIT_WIDTH_1 = 16;
defparam sdpb_inst_41.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_41.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_41.RESET_MODE = "SYNC";

SDPB sdpb_inst_42 (
    .DO({sdpb_inst_42_dout_w[15:0],sdpb_inst_42_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_42}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_106}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_42.READ_MODE = 1'b0;
defparam sdpb_inst_42.BIT_WIDTH_0 = 16;
defparam sdpb_inst_42.BIT_WIDTH_1 = 16;
defparam sdpb_inst_42.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_42.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_42.RESET_MODE = "SYNC";

SDPB sdpb_inst_43 (
    .DO({sdpb_inst_43_dout_w[15:0],sdpb_inst_43_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_43}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_107}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_43.READ_MODE = 1'b0;
defparam sdpb_inst_43.BIT_WIDTH_0 = 16;
defparam sdpb_inst_43.BIT_WIDTH_1 = 16;
defparam sdpb_inst_43.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_43.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_43.RESET_MODE = "SYNC";

SDPB sdpb_inst_44 (
    .DO({sdpb_inst_44_dout_w[15:0],sdpb_inst_44_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_44}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_108}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_44.READ_MODE = 1'b0;
defparam sdpb_inst_44.BIT_WIDTH_0 = 16;
defparam sdpb_inst_44.BIT_WIDTH_1 = 16;
defparam sdpb_inst_44.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_44.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_44.RESET_MODE = "SYNC";

SDPB sdpb_inst_45 (
    .DO({sdpb_inst_45_dout_w[15:0],sdpb_inst_45_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_45}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_109}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_45.READ_MODE = 1'b0;
defparam sdpb_inst_45.BIT_WIDTH_0 = 16;
defparam sdpb_inst_45.BIT_WIDTH_1 = 16;
defparam sdpb_inst_45.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_45.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_45.RESET_MODE = "SYNC";

SDPB sdpb_inst_46 (
    .DO({sdpb_inst_46_dout_w[15:0],sdpb_inst_46_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_46}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_110}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_46.READ_MODE = 1'b0;
defparam sdpb_inst_46.BIT_WIDTH_0 = 16;
defparam sdpb_inst_46.BIT_WIDTH_1 = 16;
defparam sdpb_inst_46.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_46.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_46.RESET_MODE = "SYNC";

SDPB sdpb_inst_47 (
    .DO({sdpb_inst_47_dout_w[15:0],sdpb_inst_47_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_47}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_111}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_47.READ_MODE = 1'b0;
defparam sdpb_inst_47.BIT_WIDTH_0 = 16;
defparam sdpb_inst_47.BIT_WIDTH_1 = 16;
defparam sdpb_inst_47.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_47.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_47.RESET_MODE = "SYNC";

SDPB sdpb_inst_48 (
    .DO({sdpb_inst_48_dout_w[15:0],sdpb_inst_48_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_48}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_112}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_48.READ_MODE = 1'b0;
defparam sdpb_inst_48.BIT_WIDTH_0 = 16;
defparam sdpb_inst_48.BIT_WIDTH_1 = 16;
defparam sdpb_inst_48.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_48.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_48.RESET_MODE = "SYNC";

SDPB sdpb_inst_49 (
    .DO({sdpb_inst_49_dout_w[15:0],sdpb_inst_49_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_49}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_113}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_49.READ_MODE = 1'b0;
defparam sdpb_inst_49.BIT_WIDTH_0 = 16;
defparam sdpb_inst_49.BIT_WIDTH_1 = 16;
defparam sdpb_inst_49.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_49.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_49.RESET_MODE = "SYNC";

SDPB sdpb_inst_50 (
    .DO({sdpb_inst_50_dout_w[15:0],sdpb_inst_50_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_50}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_114}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_50.READ_MODE = 1'b0;
defparam sdpb_inst_50.BIT_WIDTH_0 = 16;
defparam sdpb_inst_50.BIT_WIDTH_1 = 16;
defparam sdpb_inst_50.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_50.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_50.RESET_MODE = "SYNC";

SDPB sdpb_inst_51 (
    .DO({sdpb_inst_51_dout_w[15:0],sdpb_inst_51_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_51}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_51.READ_MODE = 1'b0;
defparam sdpb_inst_51.BIT_WIDTH_0 = 16;
defparam sdpb_inst_51.BIT_WIDTH_1 = 16;
defparam sdpb_inst_51.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_51.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_51.RESET_MODE = "SYNC";

SDPB sdpb_inst_52 (
    .DO({sdpb_inst_52_dout_w[15:0],sdpb_inst_52_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_52}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_116}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_52.READ_MODE = 1'b0;
defparam sdpb_inst_52.BIT_WIDTH_0 = 16;
defparam sdpb_inst_52.BIT_WIDTH_1 = 16;
defparam sdpb_inst_52.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_52.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_52.RESET_MODE = "SYNC";

SDPB sdpb_inst_53 (
    .DO({sdpb_inst_53_dout_w[15:0],sdpb_inst_53_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_53}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_117}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_53.READ_MODE = 1'b0;
defparam sdpb_inst_53.BIT_WIDTH_0 = 16;
defparam sdpb_inst_53.BIT_WIDTH_1 = 16;
defparam sdpb_inst_53.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_53.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_53.RESET_MODE = "SYNC";

SDPB sdpb_inst_54 (
    .DO({sdpb_inst_54_dout_w[15:0],sdpb_inst_54_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_54}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_118}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_54.READ_MODE = 1'b0;
defparam sdpb_inst_54.BIT_WIDTH_0 = 16;
defparam sdpb_inst_54.BIT_WIDTH_1 = 16;
defparam sdpb_inst_54.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_54.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_54.RESET_MODE = "SYNC";

SDPB sdpb_inst_55 (
    .DO({sdpb_inst_55_dout_w[15:0],sdpb_inst_55_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_55}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_119}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_55.READ_MODE = 1'b0;
defparam sdpb_inst_55.BIT_WIDTH_0 = 16;
defparam sdpb_inst_55.BIT_WIDTH_1 = 16;
defparam sdpb_inst_55.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_55.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_55.RESET_MODE = "SYNC";

SDPB sdpb_inst_56 (
    .DO({sdpb_inst_56_dout_w[15:0],sdpb_inst_56_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_120}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_56.READ_MODE = 1'b0;
defparam sdpb_inst_56.BIT_WIDTH_0 = 16;
defparam sdpb_inst_56.BIT_WIDTH_1 = 16;
defparam sdpb_inst_56.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_56.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_56.RESET_MODE = "SYNC";

SDPB sdpb_inst_57 (
    .DO({sdpb_inst_57_dout_w[15:0],sdpb_inst_57_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_121}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_57.READ_MODE = 1'b0;
defparam sdpb_inst_57.BIT_WIDTH_0 = 16;
defparam sdpb_inst_57.BIT_WIDTH_1 = 16;
defparam sdpb_inst_57.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_57.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_57.RESET_MODE = "SYNC";

SDPB sdpb_inst_58 (
    .DO({sdpb_inst_58_dout_w[15:0],sdpb_inst_58_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_58}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_122}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_58.READ_MODE = 1'b0;
defparam sdpb_inst_58.BIT_WIDTH_0 = 16;
defparam sdpb_inst_58.BIT_WIDTH_1 = 16;
defparam sdpb_inst_58.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_58.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_58.RESET_MODE = "SYNC";

SDPB sdpb_inst_59 (
    .DO({sdpb_inst_59_dout_w[15:0],sdpb_inst_59_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_59}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_123}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_59.READ_MODE = 1'b0;
defparam sdpb_inst_59.BIT_WIDTH_0 = 16;
defparam sdpb_inst_59.BIT_WIDTH_1 = 16;
defparam sdpb_inst_59.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_59.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_59.RESET_MODE = "SYNC";

SDPB sdpb_inst_60 (
    .DO({sdpb_inst_60_dout_w[15:0],sdpb_inst_60_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_60}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_124}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_60.READ_MODE = 1'b0;
defparam sdpb_inst_60.BIT_WIDTH_0 = 16;
defparam sdpb_inst_60.BIT_WIDTH_1 = 16;
defparam sdpb_inst_60.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_60.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_60.RESET_MODE = "SYNC";

SDPB sdpb_inst_61 (
    .DO({sdpb_inst_61_dout_w[15:0],sdpb_inst_61_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_61}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_125}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_61.READ_MODE = 1'b0;
defparam sdpb_inst_61.BIT_WIDTH_0 = 16;
defparam sdpb_inst_61.BIT_WIDTH_1 = 16;
defparam sdpb_inst_61.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_61.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_61.RESET_MODE = "SYNC";

SDPB sdpb_inst_62 (
    .DO({sdpb_inst_62_dout_w[15:0],sdpb_inst_62_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_62}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_126}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_62.READ_MODE = 1'b0;
defparam sdpb_inst_62.BIT_WIDTH_0 = 16;
defparam sdpb_inst_62.BIT_WIDTH_1 = 16;
defparam sdpb_inst_62.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_62.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_62.RESET_MODE = "SYNC";

SDPB sdpb_inst_63 (
    .DO({sdpb_inst_63_dout_w[15:0],sdpb_inst_63_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_63}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_127}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_63.READ_MODE = 1'b0;
defparam sdpb_inst_63.BIT_WIDTH_0 = 16;
defparam sdpb_inst_63.BIT_WIDTH_1 = 16;
defparam sdpb_inst_63.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_63.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_63.RESET_MODE = "SYNC";

SDPB sdpb_inst_64 (
    .DO({sdpb_inst_64_dout_w[15:0],sdpb_inst_64_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_64}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_64.READ_MODE = 1'b0;
defparam sdpb_inst_64.BIT_WIDTH_0 = 16;
defparam sdpb_inst_64.BIT_WIDTH_1 = 16;
defparam sdpb_inst_64.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_64.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_64.RESET_MODE = "SYNC";

SDPB sdpb_inst_65 (
    .DO({sdpb_inst_65_dout_w[15:0],sdpb_inst_65_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_65}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_65.READ_MODE = 1'b0;
defparam sdpb_inst_65.BIT_WIDTH_0 = 16;
defparam sdpb_inst_65.BIT_WIDTH_1 = 16;
defparam sdpb_inst_65.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_65.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_65.RESET_MODE = "SYNC";

SDPB sdpb_inst_66 (
    .DO({sdpb_inst_66_dout_w[15:0],sdpb_inst_66_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_66}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_66.READ_MODE = 1'b0;
defparam sdpb_inst_66.BIT_WIDTH_0 = 16;
defparam sdpb_inst_66.BIT_WIDTH_1 = 16;
defparam sdpb_inst_66.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_66.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_66.RESET_MODE = "SYNC";

SDPB sdpb_inst_67 (
    .DO({sdpb_inst_67_dout_w[15:0],sdpb_inst_67_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_67}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_67.READ_MODE = 1'b0;
defparam sdpb_inst_67.BIT_WIDTH_0 = 16;
defparam sdpb_inst_67.BIT_WIDTH_1 = 16;
defparam sdpb_inst_67.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_67.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_67.RESET_MODE = "SYNC";

SDPB sdpb_inst_68 (
    .DO({sdpb_inst_68_dout_w[15:0],sdpb_inst_68_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_68}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_68.READ_MODE = 1'b0;
defparam sdpb_inst_68.BIT_WIDTH_0 = 16;
defparam sdpb_inst_68.BIT_WIDTH_1 = 16;
defparam sdpb_inst_68.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_68.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_68.RESET_MODE = "SYNC";

SDPB sdpb_inst_69 (
    .DO({sdpb_inst_69_dout_w[15:0],sdpb_inst_69_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_69}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_69.READ_MODE = 1'b0;
defparam sdpb_inst_69.BIT_WIDTH_0 = 16;
defparam sdpb_inst_69.BIT_WIDTH_1 = 16;
defparam sdpb_inst_69.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_69.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_69.RESET_MODE = "SYNC";

SDPB sdpb_inst_70 (
    .DO({sdpb_inst_70_dout_w[15:0],sdpb_inst_70_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_70}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_70.READ_MODE = 1'b0;
defparam sdpb_inst_70.BIT_WIDTH_0 = 16;
defparam sdpb_inst_70.BIT_WIDTH_1 = 16;
defparam sdpb_inst_70.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_70.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_70.RESET_MODE = "SYNC";

SDPB sdpb_inst_71 (
    .DO({sdpb_inst_71_dout_w[15:0],sdpb_inst_71_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_71}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_71.READ_MODE = 1'b0;
defparam sdpb_inst_71.BIT_WIDTH_0 = 16;
defparam sdpb_inst_71.BIT_WIDTH_1 = 16;
defparam sdpb_inst_71.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_71.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_71.RESET_MODE = "SYNC";

SDPB sdpb_inst_72 (
    .DO({sdpb_inst_72_dout_w[15:0],sdpb_inst_72_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_72}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_72.READ_MODE = 1'b0;
defparam sdpb_inst_72.BIT_WIDTH_0 = 16;
defparam sdpb_inst_72.BIT_WIDTH_1 = 16;
defparam sdpb_inst_72.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_72.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_72.RESET_MODE = "SYNC";

SDPB sdpb_inst_73 (
    .DO({sdpb_inst_73_dout_w[15:0],sdpb_inst_73_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_73}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_73.READ_MODE = 1'b0;
defparam sdpb_inst_73.BIT_WIDTH_0 = 16;
defparam sdpb_inst_73.BIT_WIDTH_1 = 16;
defparam sdpb_inst_73.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_73.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_73.RESET_MODE = "SYNC";

SDPB sdpb_inst_74 (
    .DO({sdpb_inst_74_dout_w[15:0],sdpb_inst_74_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_74}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_74.READ_MODE = 1'b0;
defparam sdpb_inst_74.BIT_WIDTH_0 = 16;
defparam sdpb_inst_74.BIT_WIDTH_1 = 16;
defparam sdpb_inst_74.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_74.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_74.RESET_MODE = "SYNC";

SDPB sdpb_inst_75 (
    .DO({sdpb_inst_75_dout_w[15:0],sdpb_inst_75_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_75}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_75.READ_MODE = 1'b0;
defparam sdpb_inst_75.BIT_WIDTH_0 = 16;
defparam sdpb_inst_75.BIT_WIDTH_1 = 16;
defparam sdpb_inst_75.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_75.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_75.RESET_MODE = "SYNC";

SDPB sdpb_inst_76 (
    .DO({sdpb_inst_76_dout_w[15:0],sdpb_inst_76_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_76}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_76.READ_MODE = 1'b0;
defparam sdpb_inst_76.BIT_WIDTH_0 = 16;
defparam sdpb_inst_76.BIT_WIDTH_1 = 16;
defparam sdpb_inst_76.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_76.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_76.RESET_MODE = "SYNC";

SDPB sdpb_inst_77 (
    .DO({sdpb_inst_77_dout_w[15:0],sdpb_inst_77_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_77}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_77.READ_MODE = 1'b0;
defparam sdpb_inst_77.BIT_WIDTH_0 = 16;
defparam sdpb_inst_77.BIT_WIDTH_1 = 16;
defparam sdpb_inst_77.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_77.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_77.RESET_MODE = "SYNC";

SDPB sdpb_inst_78 (
    .DO({sdpb_inst_78_dout_w[15:0],sdpb_inst_78_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_78}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_78.READ_MODE = 1'b0;
defparam sdpb_inst_78.BIT_WIDTH_0 = 16;
defparam sdpb_inst_78.BIT_WIDTH_1 = 16;
defparam sdpb_inst_78.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_78.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_78.RESET_MODE = "SYNC";

SDPB sdpb_inst_79 (
    .DO({sdpb_inst_79_dout_w[15:0],sdpb_inst_79_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_79}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_79.READ_MODE = 1'b0;
defparam sdpb_inst_79.BIT_WIDTH_0 = 16;
defparam sdpb_inst_79.BIT_WIDTH_1 = 16;
defparam sdpb_inst_79.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_79.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_79.RESET_MODE = "SYNC";

SDPB sdpb_inst_80 (
    .DO({sdpb_inst_80_dout_w[15:0],sdpb_inst_80_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_16}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_80}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_80.READ_MODE = 1'b0;
defparam sdpb_inst_80.BIT_WIDTH_0 = 16;
defparam sdpb_inst_80.BIT_WIDTH_1 = 16;
defparam sdpb_inst_80.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_80.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_80.RESET_MODE = "SYNC";

SDPB sdpb_inst_81 (
    .DO({sdpb_inst_81_dout_w[15:0],sdpb_inst_81_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_17}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_81}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_81.READ_MODE = 1'b0;
defparam sdpb_inst_81.BIT_WIDTH_0 = 16;
defparam sdpb_inst_81.BIT_WIDTH_1 = 16;
defparam sdpb_inst_81.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_81.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_81.RESET_MODE = "SYNC";

SDPB sdpb_inst_82 (
    .DO({sdpb_inst_82_dout_w[15:0],sdpb_inst_82_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_18}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_82}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_82.READ_MODE = 1'b0;
defparam sdpb_inst_82.BIT_WIDTH_0 = 16;
defparam sdpb_inst_82.BIT_WIDTH_1 = 16;
defparam sdpb_inst_82.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_82.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_82.RESET_MODE = "SYNC";

SDPB sdpb_inst_83 (
    .DO({sdpb_inst_83_dout_w[15:0],sdpb_inst_83_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_19}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_83}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_83.READ_MODE = 1'b0;
defparam sdpb_inst_83.BIT_WIDTH_0 = 16;
defparam sdpb_inst_83.BIT_WIDTH_1 = 16;
defparam sdpb_inst_83.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_83.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_83.RESET_MODE = "SYNC";

SDPB sdpb_inst_84 (
    .DO({sdpb_inst_84_dout_w[15:0],sdpb_inst_84_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_20}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_84}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_84.READ_MODE = 1'b0;
defparam sdpb_inst_84.BIT_WIDTH_0 = 16;
defparam sdpb_inst_84.BIT_WIDTH_1 = 16;
defparam sdpb_inst_84.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_84.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_84.RESET_MODE = "SYNC";

SDPB sdpb_inst_85 (
    .DO({sdpb_inst_85_dout_w[15:0],sdpb_inst_85_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_21}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_85}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_85.READ_MODE = 1'b0;
defparam sdpb_inst_85.BIT_WIDTH_0 = 16;
defparam sdpb_inst_85.BIT_WIDTH_1 = 16;
defparam sdpb_inst_85.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_85.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_85.RESET_MODE = "SYNC";

SDPB sdpb_inst_86 (
    .DO({sdpb_inst_86_dout_w[15:0],sdpb_inst_86_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_22}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_86}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_86.READ_MODE = 1'b0;
defparam sdpb_inst_86.BIT_WIDTH_0 = 16;
defparam sdpb_inst_86.BIT_WIDTH_1 = 16;
defparam sdpb_inst_86.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_86.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_86.RESET_MODE = "SYNC";

SDPB sdpb_inst_87 (
    .DO({sdpb_inst_87_dout_w[15:0],sdpb_inst_87_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_23}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_87}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_87.READ_MODE = 1'b0;
defparam sdpb_inst_87.BIT_WIDTH_0 = 16;
defparam sdpb_inst_87.BIT_WIDTH_1 = 16;
defparam sdpb_inst_87.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_87.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_87.RESET_MODE = "SYNC";

SDPB sdpb_inst_88 (
    .DO({sdpb_inst_88_dout_w[15:0],sdpb_inst_88_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_24}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_88}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_88.READ_MODE = 1'b0;
defparam sdpb_inst_88.BIT_WIDTH_0 = 16;
defparam sdpb_inst_88.BIT_WIDTH_1 = 16;
defparam sdpb_inst_88.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_88.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_88.RESET_MODE = "SYNC";

SDPB sdpb_inst_89 (
    .DO({sdpb_inst_89_dout_w[15:0],sdpb_inst_89_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_25}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_89}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_89.READ_MODE = 1'b0;
defparam sdpb_inst_89.BIT_WIDTH_0 = 16;
defparam sdpb_inst_89.BIT_WIDTH_1 = 16;
defparam sdpb_inst_89.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_89.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_89.RESET_MODE = "SYNC";

SDPB sdpb_inst_90 (
    .DO({sdpb_inst_90_dout_w[15:0],sdpb_inst_90_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_26}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_90}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_90.READ_MODE = 1'b0;
defparam sdpb_inst_90.BIT_WIDTH_0 = 16;
defparam sdpb_inst_90.BIT_WIDTH_1 = 16;
defparam sdpb_inst_90.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_90.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_90.RESET_MODE = "SYNC";

SDPB sdpb_inst_91 (
    .DO({sdpb_inst_91_dout_w[15:0],sdpb_inst_91_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_27}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_91}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_91.READ_MODE = 1'b0;
defparam sdpb_inst_91.BIT_WIDTH_0 = 16;
defparam sdpb_inst_91.BIT_WIDTH_1 = 16;
defparam sdpb_inst_91.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_91.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_91.RESET_MODE = "SYNC";

SDPB sdpb_inst_92 (
    .DO({sdpb_inst_92_dout_w[15:0],sdpb_inst_92_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_28}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_92}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_92.READ_MODE = 1'b0;
defparam sdpb_inst_92.BIT_WIDTH_0 = 16;
defparam sdpb_inst_92.BIT_WIDTH_1 = 16;
defparam sdpb_inst_92.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_92.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_92.RESET_MODE = "SYNC";

SDPB sdpb_inst_93 (
    .DO({sdpb_inst_93_dout_w[15:0],sdpb_inst_93_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_29}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_93}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_93.READ_MODE = 1'b0;
defparam sdpb_inst_93.BIT_WIDTH_0 = 16;
defparam sdpb_inst_93.BIT_WIDTH_1 = 16;
defparam sdpb_inst_93.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_93.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_93.RESET_MODE = "SYNC";

SDPB sdpb_inst_94 (
    .DO({sdpb_inst_94_dout_w[15:0],sdpb_inst_94_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_30}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_94}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_94.READ_MODE = 1'b0;
defparam sdpb_inst_94.BIT_WIDTH_0 = 16;
defparam sdpb_inst_94.BIT_WIDTH_1 = 16;
defparam sdpb_inst_94.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_94.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_94.RESET_MODE = "SYNC";

SDPB sdpb_inst_95 (
    .DO({sdpb_inst_95_dout_w[15:0],sdpb_inst_95_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_31}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_95}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_95.READ_MODE = 1'b0;
defparam sdpb_inst_95.BIT_WIDTH_0 = 16;
defparam sdpb_inst_95.BIT_WIDTH_1 = 16;
defparam sdpb_inst_95.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_95.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_95.RESET_MODE = "SYNC";

SDPB sdpb_inst_96 (
    .DO({sdpb_inst_96_dout_w[15:0],sdpb_inst_96_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_32}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_96}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_96.READ_MODE = 1'b0;
defparam sdpb_inst_96.BIT_WIDTH_0 = 16;
defparam sdpb_inst_96.BIT_WIDTH_1 = 16;
defparam sdpb_inst_96.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_96.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_96.RESET_MODE = "SYNC";

SDPB sdpb_inst_97 (
    .DO({sdpb_inst_97_dout_w[15:0],sdpb_inst_97_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_33}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_97}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_97.READ_MODE = 1'b0;
defparam sdpb_inst_97.BIT_WIDTH_0 = 16;
defparam sdpb_inst_97.BIT_WIDTH_1 = 16;
defparam sdpb_inst_97.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_97.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_97.RESET_MODE = "SYNC";

SDPB sdpb_inst_98 (
    .DO({sdpb_inst_98_dout_w[15:0],sdpb_inst_98_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_34}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_98}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_98.READ_MODE = 1'b0;
defparam sdpb_inst_98.BIT_WIDTH_0 = 16;
defparam sdpb_inst_98.BIT_WIDTH_1 = 16;
defparam sdpb_inst_98.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_98.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_98.RESET_MODE = "SYNC";

SDPB sdpb_inst_99 (
    .DO({sdpb_inst_99_dout_w[15:0],sdpb_inst_99_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_35}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_99}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_99.READ_MODE = 1'b0;
defparam sdpb_inst_99.BIT_WIDTH_0 = 16;
defparam sdpb_inst_99.BIT_WIDTH_1 = 16;
defparam sdpb_inst_99.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_99.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_99.RESET_MODE = "SYNC";

SDPB sdpb_inst_100 (
    .DO({sdpb_inst_100_dout_w[15:0],sdpb_inst_100_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_36}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_100}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_100.READ_MODE = 1'b0;
defparam sdpb_inst_100.BIT_WIDTH_0 = 16;
defparam sdpb_inst_100.BIT_WIDTH_1 = 16;
defparam sdpb_inst_100.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_100.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_100.RESET_MODE = "SYNC";

SDPB sdpb_inst_101 (
    .DO({sdpb_inst_101_dout_w[15:0],sdpb_inst_101_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_37}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_101}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_101.READ_MODE = 1'b0;
defparam sdpb_inst_101.BIT_WIDTH_0 = 16;
defparam sdpb_inst_101.BIT_WIDTH_1 = 16;
defparam sdpb_inst_101.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_101.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_101.RESET_MODE = "SYNC";

SDPB sdpb_inst_102 (
    .DO({sdpb_inst_102_dout_w[15:0],sdpb_inst_102_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_38}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_102}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_102.READ_MODE = 1'b0;
defparam sdpb_inst_102.BIT_WIDTH_0 = 16;
defparam sdpb_inst_102.BIT_WIDTH_1 = 16;
defparam sdpb_inst_102.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_102.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_102.RESET_MODE = "SYNC";

SDPB sdpb_inst_103 (
    .DO({sdpb_inst_103_dout_w[15:0],sdpb_inst_103_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_39}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_103}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_103.READ_MODE = 1'b0;
defparam sdpb_inst_103.BIT_WIDTH_0 = 16;
defparam sdpb_inst_103.BIT_WIDTH_1 = 16;
defparam sdpb_inst_103.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_103.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_103.RESET_MODE = "SYNC";

SDPB sdpb_inst_104 (
    .DO({sdpb_inst_104_dout_w[15:0],sdpb_inst_104_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_40}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_104}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_104.READ_MODE = 1'b0;
defparam sdpb_inst_104.BIT_WIDTH_0 = 16;
defparam sdpb_inst_104.BIT_WIDTH_1 = 16;
defparam sdpb_inst_104.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_104.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_104.RESET_MODE = "SYNC";

SDPB sdpb_inst_105 (
    .DO({sdpb_inst_105_dout_w[15:0],sdpb_inst_105_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_41}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_105}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_105.READ_MODE = 1'b0;
defparam sdpb_inst_105.BIT_WIDTH_0 = 16;
defparam sdpb_inst_105.BIT_WIDTH_1 = 16;
defparam sdpb_inst_105.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_105.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_105.RESET_MODE = "SYNC";

SDPB sdpb_inst_106 (
    .DO({sdpb_inst_106_dout_w[15:0],sdpb_inst_106_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_42}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_106}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_106.READ_MODE = 1'b0;
defparam sdpb_inst_106.BIT_WIDTH_0 = 16;
defparam sdpb_inst_106.BIT_WIDTH_1 = 16;
defparam sdpb_inst_106.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_106.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_106.RESET_MODE = "SYNC";

SDPB sdpb_inst_107 (
    .DO({sdpb_inst_107_dout_w[15:0],sdpb_inst_107_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_43}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_107}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_107.READ_MODE = 1'b0;
defparam sdpb_inst_107.BIT_WIDTH_0 = 16;
defparam sdpb_inst_107.BIT_WIDTH_1 = 16;
defparam sdpb_inst_107.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_107.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_107.RESET_MODE = "SYNC";

SDPB sdpb_inst_108 (
    .DO({sdpb_inst_108_dout_w[15:0],sdpb_inst_108_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_44}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_108}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_108.READ_MODE = 1'b0;
defparam sdpb_inst_108.BIT_WIDTH_0 = 16;
defparam sdpb_inst_108.BIT_WIDTH_1 = 16;
defparam sdpb_inst_108.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_108.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_108.RESET_MODE = "SYNC";

SDPB sdpb_inst_109 (
    .DO({sdpb_inst_109_dout_w[15:0],sdpb_inst_109_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_45}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_109}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_109.READ_MODE = 1'b0;
defparam sdpb_inst_109.BIT_WIDTH_0 = 16;
defparam sdpb_inst_109.BIT_WIDTH_1 = 16;
defparam sdpb_inst_109.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_109.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_109.RESET_MODE = "SYNC";

SDPB sdpb_inst_110 (
    .DO({sdpb_inst_110_dout_w[15:0],sdpb_inst_110_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_46}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_110}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_110.READ_MODE = 1'b0;
defparam sdpb_inst_110.BIT_WIDTH_0 = 16;
defparam sdpb_inst_110.BIT_WIDTH_1 = 16;
defparam sdpb_inst_110.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_110.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_110.RESET_MODE = "SYNC";

SDPB sdpb_inst_111 (
    .DO({sdpb_inst_111_dout_w[15:0],sdpb_inst_111_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_47}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_111}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_111.READ_MODE = 1'b0;
defparam sdpb_inst_111.BIT_WIDTH_0 = 16;
defparam sdpb_inst_111.BIT_WIDTH_1 = 16;
defparam sdpb_inst_111.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_111.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_111.RESET_MODE = "SYNC";

SDPB sdpb_inst_112 (
    .DO({sdpb_inst_112_dout_w[15:0],sdpb_inst_112_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_48}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_112}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_112.READ_MODE = 1'b0;
defparam sdpb_inst_112.BIT_WIDTH_0 = 16;
defparam sdpb_inst_112.BIT_WIDTH_1 = 16;
defparam sdpb_inst_112.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_112.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_112.RESET_MODE = "SYNC";

SDPB sdpb_inst_113 (
    .DO({sdpb_inst_113_dout_w[15:0],sdpb_inst_113_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_49}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_113}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_113.READ_MODE = 1'b0;
defparam sdpb_inst_113.BIT_WIDTH_0 = 16;
defparam sdpb_inst_113.BIT_WIDTH_1 = 16;
defparam sdpb_inst_113.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_113.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_113.RESET_MODE = "SYNC";

SDPB sdpb_inst_114 (
    .DO({sdpb_inst_114_dout_w[15:0],sdpb_inst_114_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_50}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_114}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_114.READ_MODE = 1'b0;
defparam sdpb_inst_114.BIT_WIDTH_0 = 16;
defparam sdpb_inst_114.BIT_WIDTH_1 = 16;
defparam sdpb_inst_114.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_114.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_114.RESET_MODE = "SYNC";

SDPB sdpb_inst_115 (
    .DO({sdpb_inst_115_dout_w[15:0],sdpb_inst_115_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_51}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_115.READ_MODE = 1'b0;
defparam sdpb_inst_115.BIT_WIDTH_0 = 16;
defparam sdpb_inst_115.BIT_WIDTH_1 = 16;
defparam sdpb_inst_115.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_115.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_115.RESET_MODE = "SYNC";

SDPB sdpb_inst_116 (
    .DO({sdpb_inst_116_dout_w[15:0],sdpb_inst_116_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_52}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_116}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_116.READ_MODE = 1'b0;
defparam sdpb_inst_116.BIT_WIDTH_0 = 16;
defparam sdpb_inst_116.BIT_WIDTH_1 = 16;
defparam sdpb_inst_116.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_116.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_116.RESET_MODE = "SYNC";

SDPB sdpb_inst_117 (
    .DO({sdpb_inst_117_dout_w[15:0],sdpb_inst_117_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_53}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_117}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_117.READ_MODE = 1'b0;
defparam sdpb_inst_117.BIT_WIDTH_0 = 16;
defparam sdpb_inst_117.BIT_WIDTH_1 = 16;
defparam sdpb_inst_117.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_117.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_117.RESET_MODE = "SYNC";

SDPB sdpb_inst_118 (
    .DO({sdpb_inst_118_dout_w[15:0],sdpb_inst_118_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_54}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_118}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_118.READ_MODE = 1'b0;
defparam sdpb_inst_118.BIT_WIDTH_0 = 16;
defparam sdpb_inst_118.BIT_WIDTH_1 = 16;
defparam sdpb_inst_118.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_118.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_118.RESET_MODE = "SYNC";

SDPB sdpb_inst_119 (
    .DO({sdpb_inst_119_dout_w[15:0],sdpb_inst_119_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_55}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_119}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_119.READ_MODE = 1'b0;
defparam sdpb_inst_119.BIT_WIDTH_0 = 16;
defparam sdpb_inst_119.BIT_WIDTH_1 = 16;
defparam sdpb_inst_119.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_119.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_119.RESET_MODE = "SYNC";

SDPB sdpb_inst_120 (
    .DO({sdpb_inst_120_dout_w[15:0],sdpb_inst_120_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_120}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_120.READ_MODE = 1'b0;
defparam sdpb_inst_120.BIT_WIDTH_0 = 16;
defparam sdpb_inst_120.BIT_WIDTH_1 = 16;
defparam sdpb_inst_120.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_120.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_120.RESET_MODE = "SYNC";

SDPB sdpb_inst_121 (
    .DO({sdpb_inst_121_dout_w[15:0],sdpb_inst_121_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_121}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_121.READ_MODE = 1'b0;
defparam sdpb_inst_121.BIT_WIDTH_0 = 16;
defparam sdpb_inst_121.BIT_WIDTH_1 = 16;
defparam sdpb_inst_121.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_121.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_121.RESET_MODE = "SYNC";

SDPB sdpb_inst_122 (
    .DO({sdpb_inst_122_dout_w[15:0],sdpb_inst_122_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_58}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_122}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_122.READ_MODE = 1'b0;
defparam sdpb_inst_122.BIT_WIDTH_0 = 16;
defparam sdpb_inst_122.BIT_WIDTH_1 = 16;
defparam sdpb_inst_122.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_122.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_122.RESET_MODE = "SYNC";

SDPB sdpb_inst_123 (
    .DO({sdpb_inst_123_dout_w[15:0],sdpb_inst_123_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_59}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_123}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_123.READ_MODE = 1'b0;
defparam sdpb_inst_123.BIT_WIDTH_0 = 16;
defparam sdpb_inst_123.BIT_WIDTH_1 = 16;
defparam sdpb_inst_123.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_123.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_123.RESET_MODE = "SYNC";

SDPB sdpb_inst_124 (
    .DO({sdpb_inst_124_dout_w[15:0],sdpb_inst_124_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_60}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_124}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_124.READ_MODE = 1'b0;
defparam sdpb_inst_124.BIT_WIDTH_0 = 16;
defparam sdpb_inst_124.BIT_WIDTH_1 = 16;
defparam sdpb_inst_124.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_124.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_124.RESET_MODE = "SYNC";

SDPB sdpb_inst_125 (
    .DO({sdpb_inst_125_dout_w[15:0],sdpb_inst_125_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_61}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_125}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_125.READ_MODE = 1'b0;
defparam sdpb_inst_125.BIT_WIDTH_0 = 16;
defparam sdpb_inst_125.BIT_WIDTH_1 = 16;
defparam sdpb_inst_125.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_125.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_125.RESET_MODE = "SYNC";

SDPB sdpb_inst_126 (
    .DO({sdpb_inst_126_dout_w[15:0],sdpb_inst_126_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_62}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_126}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_126.READ_MODE = 1'b0;
defparam sdpb_inst_126.BIT_WIDTH_0 = 16;
defparam sdpb_inst_126.BIT_WIDTH_1 = 16;
defparam sdpb_inst_126.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_126.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_126.RESET_MODE = "SYNC";

SDPB sdpb_inst_127 (
    .DO({sdpb_inst_127_dout_w[15:0],sdpb_inst_127_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_63}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_127}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_127.READ_MODE = 1'b0;
defparam sdpb_inst_127.BIT_WIDTH_0 = 16;
defparam sdpb_inst_127.BIT_WIDTH_1 = 16;
defparam sdpb_inst_127.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_127.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_127.RESET_MODE = "SYNC";

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[10]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sdpb_inst_2_dout[0]),
  .I1(sdpb_inst_3_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sdpb_inst_4_dout[0]),
  .I1(sdpb_inst_5_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sdpb_inst_6_dout[0]),
  .I1(sdpb_inst_7_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sdpb_inst_8_dout[0]),
  .I1(sdpb_inst_9_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sdpb_inst_10_dout[0]),
  .I1(sdpb_inst_11_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sdpb_inst_12_dout[0]),
  .I1(sdpb_inst_13_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(sdpb_inst_14_dout[0]),
  .I1(sdpb_inst_15_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sdpb_inst_16_dout[0]),
  .I1(sdpb_inst_17_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(sdpb_inst_18_dout[0]),
  .I1(sdpb_inst_19_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(sdpb_inst_20_dout[0]),
  .I1(sdpb_inst_21_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(sdpb_inst_22_dout[0]),
  .I1(sdpb_inst_23_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(sdpb_inst_24_dout[0]),
  .I1(sdpb_inst_25_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(sdpb_inst_26_dout[0]),
  .I1(sdpb_inst_27_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(sdpb_inst_28_dout[0]),
  .I1(sdpb_inst_29_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sdpb_inst_30_dout[0]),
  .I1(sdpb_inst_31_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sdpb_inst_32_dout[0]),
  .I1(sdpb_inst_33_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(sdpb_inst_34_dout[0]),
  .I1(sdpb_inst_35_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(sdpb_inst_36_dout[0]),
  .I1(sdpb_inst_37_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(sdpb_inst_38_dout[0]),
  .I1(sdpb_inst_39_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(sdpb_inst_40_dout[0]),
  .I1(sdpb_inst_41_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sdpb_inst_42_dout[0]),
  .I1(sdpb_inst_43_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(sdpb_inst_44_dout[0]),
  .I1(sdpb_inst_45_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(sdpb_inst_46_dout[0]),
  .I1(sdpb_inst_47_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(sdpb_inst_48_dout[0]),
  .I1(sdpb_inst_49_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(sdpb_inst_50_dout[0]),
  .I1(sdpb_inst_51_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(sdpb_inst_52_dout[0]),
  .I1(sdpb_inst_53_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(sdpb_inst_54_dout[0]),
  .I1(sdpb_inst_55_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(sdpb_inst_56_dout[0]),
  .I1(sdpb_inst_57_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(sdpb_inst_58_dout[0]),
  .I1(sdpb_inst_59_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(sdpb_inst_60_dout[0]),
  .I1(sdpb_inst_61_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(sdpb_inst_62_dout[0]),
  .I1(sdpb_inst_63_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_4)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_4)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_4)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_4)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_4)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_4)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_4)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_4)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_4)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_4)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(dff_q_4)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(dff_q_4)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(dff_q_4)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(dff_q_4)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_4)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_4)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_3)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_3)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_3)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(dff_q_3)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(dff_q_3)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_48),
  .I1(mux_o_49),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_50),
  .I1(mux_o_51),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_52),
  .I1(mux_o_53),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(dff_q_2)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(dff_q_1)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(dff_q_1)
);
MUX2 mux_inst_62 (
  .O(dout[0]),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_0)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sdpb_inst_0_dout[1]),
  .I1(sdpb_inst_1_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sdpb_inst_2_dout[1]),
  .I1(sdpb_inst_3_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(sdpb_inst_4_dout[1]),
  .I1(sdpb_inst_5_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sdpb_inst_6_dout[1]),
  .I1(sdpb_inst_7_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sdpb_inst_8_dout[1]),
  .I1(sdpb_inst_9_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(sdpb_inst_10_dout[1]),
  .I1(sdpb_inst_11_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(sdpb_inst_12_dout[1]),
  .I1(sdpb_inst_13_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(sdpb_inst_14_dout[1]),
  .I1(sdpb_inst_15_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(sdpb_inst_16_dout[1]),
  .I1(sdpb_inst_17_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(sdpb_inst_18_dout[1]),
  .I1(sdpb_inst_19_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(sdpb_inst_20_dout[1]),
  .I1(sdpb_inst_21_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(sdpb_inst_22_dout[1]),
  .I1(sdpb_inst_23_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(sdpb_inst_24_dout[1]),
  .I1(sdpb_inst_25_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sdpb_inst_26_dout[1]),
  .I1(sdpb_inst_27_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(sdpb_inst_28_dout[1]),
  .I1(sdpb_inst_29_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sdpb_inst_30_dout[1]),
  .I1(sdpb_inst_31_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(sdpb_inst_32_dout[1]),
  .I1(sdpb_inst_33_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(sdpb_inst_34_dout[1]),
  .I1(sdpb_inst_35_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(sdpb_inst_36_dout[1]),
  .I1(sdpb_inst_37_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(sdpb_inst_38_dout[1]),
  .I1(sdpb_inst_39_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(sdpb_inst_40_dout[1]),
  .I1(sdpb_inst_41_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(sdpb_inst_42_dout[1]),
  .I1(sdpb_inst_43_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(sdpb_inst_44_dout[1]),
  .I1(sdpb_inst_45_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(sdpb_inst_46_dout[1]),
  .I1(sdpb_inst_47_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(sdpb_inst_48_dout[1]),
  .I1(sdpb_inst_49_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(sdpb_inst_50_dout[1]),
  .I1(sdpb_inst_51_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(sdpb_inst_52_dout[1]),
  .I1(sdpb_inst_53_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(sdpb_inst_54_dout[1]),
  .I1(sdpb_inst_55_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(sdpb_inst_56_dout[1]),
  .I1(sdpb_inst_57_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(sdpb_inst_58_dout[1]),
  .I1(sdpb_inst_59_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(sdpb_inst_60_dout[1]),
  .I1(sdpb_inst_61_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(sdpb_inst_62_dout[1]),
  .I1(sdpb_inst_63_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_63),
  .I1(mux_o_64),
  .S0(dff_q_4)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_65),
  .I1(mux_o_66),
  .S0(dff_q_4)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_67),
  .I1(mux_o_68),
  .S0(dff_q_4)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_69),
  .I1(mux_o_70),
  .S0(dff_q_4)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_71),
  .I1(mux_o_72),
  .S0(dff_q_4)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_73),
  .I1(mux_o_74),
  .S0(dff_q_4)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(dff_q_4)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_4)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_4)
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_4)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_4)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_4)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(dff_q_4)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(mux_o_89),
  .I1(mux_o_90),
  .S0(dff_q_4)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_91),
  .I1(mux_o_92),
  .S0(dff_q_4)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(dff_q_4)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_99),
  .I1(mux_o_100),
  .S0(dff_q_3)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(dff_q_3)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_103),
  .I1(mux_o_104),
  .S0(dff_q_3)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_3)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_3)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_3)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(dff_q_2)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_2)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(dff_q_1)
);
MUX2 mux_inst_125 (
  .O(dout[1]),
  .I0(mux_o_123),
  .I1(mux_o_124),
  .S0(dff_q_0)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(sdpb_inst_0_dout[2]),
  .I1(sdpb_inst_1_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(sdpb_inst_2_dout[2]),
  .I1(sdpb_inst_3_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(sdpb_inst_4_dout[2]),
  .I1(sdpb_inst_5_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(sdpb_inst_6_dout[2]),
  .I1(sdpb_inst_7_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(sdpb_inst_8_dout[2]),
  .I1(sdpb_inst_9_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(sdpb_inst_10_dout[2]),
  .I1(sdpb_inst_11_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(sdpb_inst_12_dout[2]),
  .I1(sdpb_inst_13_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(sdpb_inst_14_dout[2]),
  .I1(sdpb_inst_15_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(sdpb_inst_16_dout[2]),
  .I1(sdpb_inst_17_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(sdpb_inst_18_dout[2]),
  .I1(sdpb_inst_19_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sdpb_inst_20_dout[2]),
  .I1(sdpb_inst_21_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(sdpb_inst_22_dout[2]),
  .I1(sdpb_inst_23_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(sdpb_inst_24_dout[2]),
  .I1(sdpb_inst_25_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(sdpb_inst_26_dout[2]),
  .I1(sdpb_inst_27_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(sdpb_inst_28_dout[2]),
  .I1(sdpb_inst_29_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(sdpb_inst_30_dout[2]),
  .I1(sdpb_inst_31_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(sdpb_inst_32_dout[2]),
  .I1(sdpb_inst_33_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(sdpb_inst_34_dout[2]),
  .I1(sdpb_inst_35_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(sdpb_inst_36_dout[2]),
  .I1(sdpb_inst_37_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(sdpb_inst_38_dout[2]),
  .I1(sdpb_inst_39_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(sdpb_inst_40_dout[2]),
  .I1(sdpb_inst_41_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(sdpb_inst_42_dout[2]),
  .I1(sdpb_inst_43_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(sdpb_inst_44_dout[2]),
  .I1(sdpb_inst_45_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(sdpb_inst_46_dout[2]),
  .I1(sdpb_inst_47_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(sdpb_inst_48_dout[2]),
  .I1(sdpb_inst_49_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(sdpb_inst_50_dout[2]),
  .I1(sdpb_inst_51_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(sdpb_inst_52_dout[2]),
  .I1(sdpb_inst_53_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(sdpb_inst_54_dout[2]),
  .I1(sdpb_inst_55_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(sdpb_inst_56_dout[2]),
  .I1(sdpb_inst_57_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(sdpb_inst_58_dout[2]),
  .I1(sdpb_inst_59_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(sdpb_inst_60_dout[2]),
  .I1(sdpb_inst_61_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(sdpb_inst_62_dout[2]),
  .I1(sdpb_inst_63_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_4)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_4)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_4)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(dff_q_4)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_134),
  .I1(mux_o_135),
  .S0(dff_q_4)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_136),
  .I1(mux_o_137),
  .S0(dff_q_4)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(mux_o_138),
  .I1(mux_o_139),
  .S0(dff_q_4)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(dff_q_4)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_4)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_4)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_4)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(dff_q_4)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_4)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_4)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_4)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_4)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_3)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(dff_q_3)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(dff_q_3)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_164),
  .I1(mux_o_165),
  .S0(dff_q_3)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_166),
  .I1(mux_o_167),
  .S0(dff_q_3)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(dff_q_3)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(dff_q_3)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(dff_q_3)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(mux_o_174),
  .I1(mux_o_175),
  .S0(dff_q_2)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_176),
  .I1(mux_o_177),
  .S0(dff_q_2)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_178),
  .I1(mux_o_179),
  .S0(dff_q_2)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(dff_q_2)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_1)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_1)
);
MUX2 mux_inst_188 (
  .O(dout[2]),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_0)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(sdpb_inst_0_dout[3]),
  .I1(sdpb_inst_1_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(sdpb_inst_2_dout[3]),
  .I1(sdpb_inst_3_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(sdpb_inst_4_dout[3]),
  .I1(sdpb_inst_5_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(sdpb_inst_6_dout[3]),
  .I1(sdpb_inst_7_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(sdpb_inst_8_dout[3]),
  .I1(sdpb_inst_9_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(sdpb_inst_10_dout[3]),
  .I1(sdpb_inst_11_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(sdpb_inst_12_dout[3]),
  .I1(sdpb_inst_13_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(sdpb_inst_14_dout[3]),
  .I1(sdpb_inst_15_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sdpb_inst_16_dout[3]),
  .I1(sdpb_inst_17_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(sdpb_inst_18_dout[3]),
  .I1(sdpb_inst_19_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(sdpb_inst_20_dout[3]),
  .I1(sdpb_inst_21_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(sdpb_inst_22_dout[3]),
  .I1(sdpb_inst_23_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(sdpb_inst_24_dout[3]),
  .I1(sdpb_inst_25_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(sdpb_inst_26_dout[3]),
  .I1(sdpb_inst_27_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(sdpb_inst_28_dout[3]),
  .I1(sdpb_inst_29_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(sdpb_inst_30_dout[3]),
  .I1(sdpb_inst_31_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(sdpb_inst_32_dout[3]),
  .I1(sdpb_inst_33_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(sdpb_inst_34_dout[3]),
  .I1(sdpb_inst_35_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(sdpb_inst_36_dout[3]),
  .I1(sdpb_inst_37_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(sdpb_inst_38_dout[3]),
  .I1(sdpb_inst_39_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(sdpb_inst_40_dout[3]),
  .I1(sdpb_inst_41_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(sdpb_inst_42_dout[3]),
  .I1(sdpb_inst_43_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(sdpb_inst_44_dout[3]),
  .I1(sdpb_inst_45_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(sdpb_inst_46_dout[3]),
  .I1(sdpb_inst_47_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(sdpb_inst_48_dout[3]),
  .I1(sdpb_inst_49_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(sdpb_inst_50_dout[3]),
  .I1(sdpb_inst_51_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(sdpb_inst_52_dout[3]),
  .I1(sdpb_inst_53_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(sdpb_inst_54_dout[3]),
  .I1(sdpb_inst_55_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(sdpb_inst_56_dout[3]),
  .I1(sdpb_inst_57_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(sdpb_inst_58_dout[3]),
  .I1(sdpb_inst_59_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(sdpb_inst_60_dout[3]),
  .I1(sdpb_inst_61_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(sdpb_inst_62_dout[3]),
  .I1(sdpb_inst_63_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_4)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(dff_q_4)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(dff_q_4)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(dff_q_4)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(dff_q_4)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(dff_q_4)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_4)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_4)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_4)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_4)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(mux_o_209),
  .I1(mux_o_210),
  .S0(dff_q_4)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(mux_o_211),
  .I1(mux_o_212),
  .S0(dff_q_4)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_213),
  .I1(mux_o_214),
  .S0(dff_q_4)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_215),
  .I1(mux_o_216),
  .S0(dff_q_4)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_4)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_4)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_3)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(dff_q_3)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_3)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_3)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_3)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_3)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_2)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_2)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(dff_q_2)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(dff_q_2)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_1)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_247),
  .I1(mux_o_248),
  .S0(dff_q_1)
);
MUX2 mux_inst_251 (
  .O(dout[3]),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(dff_q_0)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(sdpb_inst_0_dout[4]),
  .I1(sdpb_inst_1_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(sdpb_inst_2_dout[4]),
  .I1(sdpb_inst_3_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(sdpb_inst_4_dout[4]),
  .I1(sdpb_inst_5_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(sdpb_inst_6_dout[4]),
  .I1(sdpb_inst_7_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(sdpb_inst_8_dout[4]),
  .I1(sdpb_inst_9_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(sdpb_inst_10_dout[4]),
  .I1(sdpb_inst_11_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(sdpb_inst_12_dout[4]),
  .I1(sdpb_inst_13_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(sdpb_inst_14_dout[4]),
  .I1(sdpb_inst_15_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(sdpb_inst_16_dout[4]),
  .I1(sdpb_inst_17_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sdpb_inst_18_dout[4]),
  .I1(sdpb_inst_19_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(sdpb_inst_20_dout[4]),
  .I1(sdpb_inst_21_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(sdpb_inst_22_dout[4]),
  .I1(sdpb_inst_23_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(sdpb_inst_24_dout[4]),
  .I1(sdpb_inst_25_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(sdpb_inst_26_dout[4]),
  .I1(sdpb_inst_27_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(sdpb_inst_28_dout[4]),
  .I1(sdpb_inst_29_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(sdpb_inst_30_dout[4]),
  .I1(sdpb_inst_31_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(sdpb_inst_32_dout[4]),
  .I1(sdpb_inst_33_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(sdpb_inst_34_dout[4]),
  .I1(sdpb_inst_35_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(sdpb_inst_36_dout[4]),
  .I1(sdpb_inst_37_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(sdpb_inst_38_dout[4]),
  .I1(sdpb_inst_39_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(sdpb_inst_40_dout[4]),
  .I1(sdpb_inst_41_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(sdpb_inst_42_dout[4]),
  .I1(sdpb_inst_43_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(sdpb_inst_44_dout[4]),
  .I1(sdpb_inst_45_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(sdpb_inst_46_dout[4]),
  .I1(sdpb_inst_47_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(sdpb_inst_48_dout[4]),
  .I1(sdpb_inst_49_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(sdpb_inst_50_dout[4]),
  .I1(sdpb_inst_51_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(sdpb_inst_52_dout[4]),
  .I1(sdpb_inst_53_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(sdpb_inst_54_dout[4]),
  .I1(sdpb_inst_55_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(sdpb_inst_56_dout[4]),
  .I1(sdpb_inst_57_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(sdpb_inst_58_dout[4]),
  .I1(sdpb_inst_59_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(sdpb_inst_60_dout[4]),
  .I1(sdpb_inst_61_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(sdpb_inst_62_dout[4]),
  .I1(sdpb_inst_63_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_4)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_4)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_4)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(dff_q_4)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(dff_q_4)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(dff_q_4)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(dff_q_4)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_4)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_4)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_4)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_4)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_4)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_4)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(dff_q_4)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_4)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_4)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_286),
  .I1(mux_o_287),
  .S0(dff_q_3)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_288),
  .I1(mux_o_289),
  .S0(dff_q_3)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_290),
  .I1(mux_o_291),
  .S0(dff_q_3)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(mux_o_292),
  .I1(mux_o_293),
  .S0(dff_q_3)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(dff_q_3)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(dff_q_3)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_3)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_2)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_2)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(dff_q_2)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(dff_q_2)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_1)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_1)
);
MUX2 mux_inst_314 (
  .O(dout[4]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_0)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sdpb_inst_0_dout[5]),
  .I1(sdpb_inst_1_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sdpb_inst_2_dout[5]),
  .I1(sdpb_inst_3_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sdpb_inst_4_dout[5]),
  .I1(sdpb_inst_5_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(sdpb_inst_6_dout[5]),
  .I1(sdpb_inst_7_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(sdpb_inst_8_dout[5]),
  .I1(sdpb_inst_9_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sdpb_inst_10_dout[5]),
  .I1(sdpb_inst_11_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sdpb_inst_12_dout[5]),
  .I1(sdpb_inst_13_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(sdpb_inst_14_dout[5]),
  .I1(sdpb_inst_15_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(sdpb_inst_16_dout[5]),
  .I1(sdpb_inst_17_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(sdpb_inst_18_dout[5]),
  .I1(sdpb_inst_19_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(sdpb_inst_20_dout[5]),
  .I1(sdpb_inst_21_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(sdpb_inst_22_dout[5]),
  .I1(sdpb_inst_23_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(sdpb_inst_24_dout[5]),
  .I1(sdpb_inst_25_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(sdpb_inst_26_dout[5]),
  .I1(sdpb_inst_27_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(sdpb_inst_28_dout[5]),
  .I1(sdpb_inst_29_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(sdpb_inst_30_dout[5]),
  .I1(sdpb_inst_31_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(sdpb_inst_32_dout[5]),
  .I1(sdpb_inst_33_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(sdpb_inst_34_dout[5]),
  .I1(sdpb_inst_35_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(sdpb_inst_36_dout[5]),
  .I1(sdpb_inst_37_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(sdpb_inst_38_dout[5]),
  .I1(sdpb_inst_39_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(sdpb_inst_40_dout[5]),
  .I1(sdpb_inst_41_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(sdpb_inst_42_dout[5]),
  .I1(sdpb_inst_43_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(sdpb_inst_44_dout[5]),
  .I1(sdpb_inst_45_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(sdpb_inst_46_dout[5]),
  .I1(sdpb_inst_47_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(sdpb_inst_48_dout[5]),
  .I1(sdpb_inst_49_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(sdpb_inst_50_dout[5]),
  .I1(sdpb_inst_51_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(sdpb_inst_52_dout[5]),
  .I1(sdpb_inst_53_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(sdpb_inst_54_dout[5]),
  .I1(sdpb_inst_55_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(sdpb_inst_56_dout[5]),
  .I1(sdpb_inst_57_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(sdpb_inst_58_dout[5]),
  .I1(sdpb_inst_59_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(sdpb_inst_60_dout[5]),
  .I1(sdpb_inst_61_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(sdpb_inst_62_dout[5]),
  .I1(sdpb_inst_63_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_4)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_4)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_4)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_321),
  .I1(mux_o_322),
  .S0(dff_q_4)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_323),
  .I1(mux_o_324),
  .S0(dff_q_4)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_325),
  .I1(mux_o_326),
  .S0(dff_q_4)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_327),
  .I1(mux_o_328),
  .S0(dff_q_4)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_329),
  .I1(mux_o_330),
  .S0(dff_q_4)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_331),
  .I1(mux_o_332),
  .S0(dff_q_4)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_333),
  .I1(mux_o_334),
  .S0(dff_q_4)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_335),
  .I1(mux_o_336),
  .S0(dff_q_4)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_337),
  .I1(mux_o_338),
  .S0(dff_q_4)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_339),
  .I1(mux_o_340),
  .S0(dff_q_4)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(dff_q_4)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_4)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_4)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(dff_q_3)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(dff_q_3)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(dff_q_3)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_3)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_359),
  .I1(mux_o_360),
  .S0(dff_q_3)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_3)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_363),
  .I1(mux_o_364),
  .S0(dff_q_2)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_365),
  .I1(mux_o_366),
  .S0(dff_q_2)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_367),
  .I1(mux_o_368),
  .S0(dff_q_2)
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(mux_o_369),
  .I1(mux_o_370),
  .S0(dff_q_2)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_371),
  .I1(mux_o_372),
  .S0(dff_q_1)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_373),
  .I1(mux_o_374),
  .S0(dff_q_1)
);
MUX2 mux_inst_377 (
  .O(dout[5]),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_0)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(sdpb_inst_0_dout[6]),
  .I1(sdpb_inst_1_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(sdpb_inst_2_dout[6]),
  .I1(sdpb_inst_3_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(sdpb_inst_4_dout[6]),
  .I1(sdpb_inst_5_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(sdpb_inst_6_dout[6]),
  .I1(sdpb_inst_7_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(sdpb_inst_8_dout[6]),
  .I1(sdpb_inst_9_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(sdpb_inst_10_dout[6]),
  .I1(sdpb_inst_11_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(sdpb_inst_12_dout[6]),
  .I1(sdpb_inst_13_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(sdpb_inst_14_dout[6]),
  .I1(sdpb_inst_15_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(sdpb_inst_16_dout[6]),
  .I1(sdpb_inst_17_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(sdpb_inst_18_dout[6]),
  .I1(sdpb_inst_19_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(sdpb_inst_20_dout[6]),
  .I1(sdpb_inst_21_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(sdpb_inst_22_dout[6]),
  .I1(sdpb_inst_23_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(sdpb_inst_24_dout[6]),
  .I1(sdpb_inst_25_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(sdpb_inst_26_dout[6]),
  .I1(sdpb_inst_27_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(sdpb_inst_28_dout[6]),
  .I1(sdpb_inst_29_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(sdpb_inst_30_dout[6]),
  .I1(sdpb_inst_31_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(sdpb_inst_32_dout[6]),
  .I1(sdpb_inst_33_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(sdpb_inst_34_dout[6]),
  .I1(sdpb_inst_35_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(sdpb_inst_36_dout[6]),
  .I1(sdpb_inst_37_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(sdpb_inst_38_dout[6]),
  .I1(sdpb_inst_39_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(sdpb_inst_40_dout[6]),
  .I1(sdpb_inst_41_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(sdpb_inst_42_dout[6]),
  .I1(sdpb_inst_43_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(sdpb_inst_44_dout[6]),
  .I1(sdpb_inst_45_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(sdpb_inst_46_dout[6]),
  .I1(sdpb_inst_47_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(sdpb_inst_48_dout[6]),
  .I1(sdpb_inst_49_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(sdpb_inst_50_dout[6]),
  .I1(sdpb_inst_51_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(sdpb_inst_52_dout[6]),
  .I1(sdpb_inst_53_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(sdpb_inst_54_dout[6]),
  .I1(sdpb_inst_55_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(sdpb_inst_56_dout[6]),
  .I1(sdpb_inst_57_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(sdpb_inst_58_dout[6]),
  .I1(sdpb_inst_59_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(sdpb_inst_60_dout[6]),
  .I1(sdpb_inst_61_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(sdpb_inst_62_dout[6]),
  .I1(sdpb_inst_63_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(dff_q_4)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(dff_q_4)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(dff_q_4)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_384),
  .I1(mux_o_385),
  .S0(dff_q_4)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_386),
  .I1(mux_o_387),
  .S0(dff_q_4)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(mux_o_388),
  .I1(mux_o_389),
  .S0(dff_q_4)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(dff_q_4)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_4)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_4)
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_4)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(dff_q_4)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(dff_q_4)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(dff_q_4)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(mux_o_404),
  .I1(mux_o_405),
  .S0(dff_q_4)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(dff_q_4)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(mux_o_408),
  .I1(mux_o_409),
  .S0(dff_q_4)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(mux_o_410),
  .I1(mux_o_411),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(mux_o_412),
  .I1(mux_o_413),
  .S0(dff_q_3)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_414),
  .I1(mux_o_415),
  .S0(dff_q_3)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_416),
  .I1(mux_o_417),
  .S0(dff_q_3)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_418),
  .I1(mux_o_419),
  .S0(dff_q_3)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(dff_q_3)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(dff_q_3)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(dff_q_3)
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(dff_q_2)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(dff_q_2)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(dff_q_2)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(dff_q_2)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(dff_q_1)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(dff_q_1)
);
MUX2 mux_inst_440 (
  .O(dout[6]),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(dff_q_0)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sdpb_inst_0_dout[7]),
  .I1(sdpb_inst_1_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sdpb_inst_2_dout[7]),
  .I1(sdpb_inst_3_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(sdpb_inst_4_dout[7]),
  .I1(sdpb_inst_5_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(sdpb_inst_6_dout[7]),
  .I1(sdpb_inst_7_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(sdpb_inst_8_dout[7]),
  .I1(sdpb_inst_9_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(sdpb_inst_10_dout[7]),
  .I1(sdpb_inst_11_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(sdpb_inst_12_dout[7]),
  .I1(sdpb_inst_13_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(sdpb_inst_14_dout[7]),
  .I1(sdpb_inst_15_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(sdpb_inst_16_dout[7]),
  .I1(sdpb_inst_17_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(sdpb_inst_18_dout[7]),
  .I1(sdpb_inst_19_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(sdpb_inst_20_dout[7]),
  .I1(sdpb_inst_21_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(sdpb_inst_22_dout[7]),
  .I1(sdpb_inst_23_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(sdpb_inst_24_dout[7]),
  .I1(sdpb_inst_25_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(sdpb_inst_26_dout[7]),
  .I1(sdpb_inst_27_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(sdpb_inst_28_dout[7]),
  .I1(sdpb_inst_29_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(sdpb_inst_30_dout[7]),
  .I1(sdpb_inst_31_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(sdpb_inst_32_dout[7]),
  .I1(sdpb_inst_33_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(sdpb_inst_34_dout[7]),
  .I1(sdpb_inst_35_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(sdpb_inst_36_dout[7]),
  .I1(sdpb_inst_37_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(sdpb_inst_38_dout[7]),
  .I1(sdpb_inst_39_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(sdpb_inst_40_dout[7]),
  .I1(sdpb_inst_41_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(sdpb_inst_42_dout[7]),
  .I1(sdpb_inst_43_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(sdpb_inst_44_dout[7]),
  .I1(sdpb_inst_45_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(sdpb_inst_46_dout[7]),
  .I1(sdpb_inst_47_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(sdpb_inst_48_dout[7]),
  .I1(sdpb_inst_49_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(sdpb_inst_50_dout[7]),
  .I1(sdpb_inst_51_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(sdpb_inst_52_dout[7]),
  .I1(sdpb_inst_53_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(sdpb_inst_54_dout[7]),
  .I1(sdpb_inst_55_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(sdpb_inst_56_dout[7]),
  .I1(sdpb_inst_57_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(sdpb_inst_58_dout[7]),
  .I1(sdpb_inst_59_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(sdpb_inst_60_dout[7]),
  .I1(sdpb_inst_61_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(sdpb_inst_62_dout[7]),
  .I1(sdpb_inst_63_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_4)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_4)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_4)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_4)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(dff_q_4)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(dff_q_4)
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(mux_o_453),
  .I1(mux_o_454),
  .S0(dff_q_4)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(mux_o_455),
  .I1(mux_o_456),
  .S0(dff_q_4)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_457),
  .I1(mux_o_458),
  .S0(dff_q_4)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_459),
  .I1(mux_o_460),
  .S0(dff_q_4)
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(dff_q_4)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_463),
  .I1(mux_o_464),
  .S0(dff_q_4)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_4)
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_4)
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_4)
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_4)
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_3)
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_3)
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_3)
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(dff_q_3)
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(dff_q_3)
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_483),
  .I1(mux_o_484),
  .S0(dff_q_3)
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(mux_o_485),
  .I1(mux_o_486),
  .S0(dff_q_3)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(mux_o_487),
  .I1(mux_o_488),
  .S0(dff_q_3)
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(mux_o_489),
  .I1(mux_o_490),
  .S0(dff_q_2)
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(dff_q_2)
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(dff_q_2)
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(mux_o_495),
  .I1(mux_o_496),
  .S0(dff_q_2)
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(mux_o_497),
  .I1(mux_o_498),
  .S0(dff_q_1)
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(mux_o_499),
  .I1(mux_o_500),
  .S0(dff_q_1)
);
MUX2 mux_inst_503 (
  .O(dout[7]),
  .I0(mux_o_501),
  .I1(mux_o_502),
  .S0(dff_q_0)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(sdpb_inst_0_dout[8]),
  .I1(sdpb_inst_1_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(sdpb_inst_2_dout[8]),
  .I1(sdpb_inst_3_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(sdpb_inst_4_dout[8]),
  .I1(sdpb_inst_5_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(sdpb_inst_6_dout[8]),
  .I1(sdpb_inst_7_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(sdpb_inst_8_dout[8]),
  .I1(sdpb_inst_9_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(sdpb_inst_10_dout[8]),
  .I1(sdpb_inst_11_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(sdpb_inst_12_dout[8]),
  .I1(sdpb_inst_13_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(sdpb_inst_14_dout[8]),
  .I1(sdpb_inst_15_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(sdpb_inst_16_dout[8]),
  .I1(sdpb_inst_17_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(sdpb_inst_18_dout[8]),
  .I1(sdpb_inst_19_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(sdpb_inst_20_dout[8]),
  .I1(sdpb_inst_21_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(sdpb_inst_22_dout[8]),
  .I1(sdpb_inst_23_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(sdpb_inst_24_dout[8]),
  .I1(sdpb_inst_25_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(sdpb_inst_26_dout[8]),
  .I1(sdpb_inst_27_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(sdpb_inst_28_dout[8]),
  .I1(sdpb_inst_29_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(sdpb_inst_30_dout[8]),
  .I1(sdpb_inst_31_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(sdpb_inst_32_dout[8]),
  .I1(sdpb_inst_33_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(sdpb_inst_34_dout[8]),
  .I1(sdpb_inst_35_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(sdpb_inst_36_dout[8]),
  .I1(sdpb_inst_37_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(sdpb_inst_38_dout[8]),
  .I1(sdpb_inst_39_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(sdpb_inst_40_dout[8]),
  .I1(sdpb_inst_41_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(sdpb_inst_42_dout[8]),
  .I1(sdpb_inst_43_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(sdpb_inst_44_dout[8]),
  .I1(sdpb_inst_45_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(sdpb_inst_46_dout[8]),
  .I1(sdpb_inst_47_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(sdpb_inst_48_dout[8]),
  .I1(sdpb_inst_49_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(sdpb_inst_50_dout[8]),
  .I1(sdpb_inst_51_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(sdpb_inst_52_dout[8]),
  .I1(sdpb_inst_53_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(sdpb_inst_54_dout[8]),
  .I1(sdpb_inst_55_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(sdpb_inst_56_dout[8]),
  .I1(sdpb_inst_57_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(sdpb_inst_58_dout[8]),
  .I1(sdpb_inst_59_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(sdpb_inst_60_dout[8]),
  .I1(sdpb_inst_61_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(sdpb_inst_62_dout[8]),
  .I1(sdpb_inst_63_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(mux_o_504),
  .I1(mux_o_505),
  .S0(dff_q_4)
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(mux_o_506),
  .I1(mux_o_507),
  .S0(dff_q_4)
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(dff_q_4)
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(dff_q_4)
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(dff_q_4)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(dff_q_4)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(dff_q_4)
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(dff_q_4)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(dff_q_4)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_4)
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(dff_q_4)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(mux_o_526),
  .I1(mux_o_527),
  .S0(dff_q_4)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(mux_o_528),
  .I1(mux_o_529),
  .S0(dff_q_4)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(mux_o_530),
  .I1(mux_o_531),
  .S0(dff_q_4)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(mux_o_532),
  .I1(mux_o_533),
  .S0(dff_q_4)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(mux_o_534),
  .I1(mux_o_535),
  .S0(dff_q_4)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(mux_o_536),
  .I1(mux_o_537),
  .S0(dff_q_3)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(mux_o_538),
  .I1(mux_o_539),
  .S0(dff_q_3)
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(dff_q_3)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(mux_o_542),
  .I1(mux_o_543),
  .S0(dff_q_3)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(dff_q_3)
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(mux_o_546),
  .I1(mux_o_547),
  .S0(dff_q_3)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(mux_o_548),
  .I1(mux_o_549),
  .S0(dff_q_3)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(mux_o_550),
  .I1(mux_o_551),
  .S0(dff_q_3)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(mux_o_552),
  .I1(mux_o_553),
  .S0(dff_q_2)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(mux_o_554),
  .I1(mux_o_555),
  .S0(dff_q_2)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(mux_o_556),
  .I1(mux_o_557),
  .S0(dff_q_2)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(dff_q_2)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(dff_q_1)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(dff_q_1)
);
MUX2 mux_inst_566 (
  .O(dout[8]),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(dff_q_0)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(sdpb_inst_0_dout[9]),
  .I1(sdpb_inst_1_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(sdpb_inst_2_dout[9]),
  .I1(sdpb_inst_3_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(sdpb_inst_4_dout[9]),
  .I1(sdpb_inst_5_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(sdpb_inst_6_dout[9]),
  .I1(sdpb_inst_7_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(sdpb_inst_8_dout[9]),
  .I1(sdpb_inst_9_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(sdpb_inst_10_dout[9]),
  .I1(sdpb_inst_11_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(sdpb_inst_12_dout[9]),
  .I1(sdpb_inst_13_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(sdpb_inst_14_dout[9]),
  .I1(sdpb_inst_15_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(sdpb_inst_16_dout[9]),
  .I1(sdpb_inst_17_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(sdpb_inst_18_dout[9]),
  .I1(sdpb_inst_19_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(sdpb_inst_20_dout[9]),
  .I1(sdpb_inst_21_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(sdpb_inst_22_dout[9]),
  .I1(sdpb_inst_23_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(sdpb_inst_24_dout[9]),
  .I1(sdpb_inst_25_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(sdpb_inst_26_dout[9]),
  .I1(sdpb_inst_27_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(sdpb_inst_28_dout[9]),
  .I1(sdpb_inst_29_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(sdpb_inst_30_dout[9]),
  .I1(sdpb_inst_31_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(sdpb_inst_32_dout[9]),
  .I1(sdpb_inst_33_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(sdpb_inst_34_dout[9]),
  .I1(sdpb_inst_35_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(sdpb_inst_36_dout[9]),
  .I1(sdpb_inst_37_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(sdpb_inst_38_dout[9]),
  .I1(sdpb_inst_39_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(sdpb_inst_40_dout[9]),
  .I1(sdpb_inst_41_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_588 (
  .O(mux_o_588),
  .I0(sdpb_inst_42_dout[9]),
  .I1(sdpb_inst_43_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(sdpb_inst_44_dout[9]),
  .I1(sdpb_inst_45_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(sdpb_inst_46_dout[9]),
  .I1(sdpb_inst_47_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(sdpb_inst_48_dout[9]),
  .I1(sdpb_inst_49_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(sdpb_inst_50_dout[9]),
  .I1(sdpb_inst_51_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(sdpb_inst_52_dout[9]),
  .I1(sdpb_inst_53_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(sdpb_inst_54_dout[9]),
  .I1(sdpb_inst_55_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(sdpb_inst_56_dout[9]),
  .I1(sdpb_inst_57_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(sdpb_inst_58_dout[9]),
  .I1(sdpb_inst_59_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(sdpb_inst_60_dout[9]),
  .I1(sdpb_inst_61_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(sdpb_inst_62_dout[9]),
  .I1(sdpb_inst_63_dout[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(mux_o_567),
  .I1(mux_o_568),
  .S0(dff_q_4)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_569),
  .I1(mux_o_570),
  .S0(dff_q_4)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_571),
  .I1(mux_o_572),
  .S0(dff_q_4)
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(mux_o_573),
  .I1(mux_o_574),
  .S0(dff_q_4)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(mux_o_575),
  .I1(mux_o_576),
  .S0(dff_q_4)
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(mux_o_577),
  .I1(mux_o_578),
  .S0(dff_q_4)
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_579),
  .I1(mux_o_580),
  .S0(dff_q_4)
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_581),
  .I1(mux_o_582),
  .S0(dff_q_4)
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_583),
  .I1(mux_o_584),
  .S0(dff_q_4)
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_585),
  .I1(mux_o_586),
  .S0(dff_q_4)
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_587),
  .I1(mux_o_588),
  .S0(dff_q_4)
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_589),
  .I1(mux_o_590),
  .S0(dff_q_4)
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_591),
  .I1(mux_o_592),
  .S0(dff_q_4)
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_593),
  .I1(mux_o_594),
  .S0(dff_q_4)
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_595),
  .I1(mux_o_596),
  .S0(dff_q_4)
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_597),
  .I1(mux_o_598),
  .S0(dff_q_4)
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_599),
  .I1(mux_o_600),
  .S0(dff_q_3)
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_601),
  .I1(mux_o_602),
  .S0(dff_q_3)
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_603),
  .I1(mux_o_604),
  .S0(dff_q_3)
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_605),
  .I1(mux_o_606),
  .S0(dff_q_3)
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(mux_o_607),
  .I1(mux_o_608),
  .S0(dff_q_3)
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(mux_o_609),
  .I1(mux_o_610),
  .S0(dff_q_3)
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(mux_o_611),
  .I1(mux_o_612),
  .S0(dff_q_3)
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(mux_o_613),
  .I1(mux_o_614),
  .S0(dff_q_3)
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(mux_o_615),
  .I1(mux_o_616),
  .S0(dff_q_2)
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_617),
  .I1(mux_o_618),
  .S0(dff_q_2)
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_619),
  .I1(mux_o_620),
  .S0(dff_q_2)
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_621),
  .I1(mux_o_622),
  .S0(dff_q_2)
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(mux_o_623),
  .I1(mux_o_624),
  .S0(dff_q_1)
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_625),
  .I1(mux_o_626),
  .S0(dff_q_1)
);
MUX2 mux_inst_629 (
  .O(dout[9]),
  .I0(mux_o_627),
  .I1(mux_o_628),
  .S0(dff_q_0)
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(sdpb_inst_0_dout[10]),
  .I1(sdpb_inst_1_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(sdpb_inst_2_dout[10]),
  .I1(sdpb_inst_3_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(sdpb_inst_4_dout[10]),
  .I1(sdpb_inst_5_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(sdpb_inst_6_dout[10]),
  .I1(sdpb_inst_7_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(sdpb_inst_8_dout[10]),
  .I1(sdpb_inst_9_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(sdpb_inst_10_dout[10]),
  .I1(sdpb_inst_11_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(sdpb_inst_12_dout[10]),
  .I1(sdpb_inst_13_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(sdpb_inst_14_dout[10]),
  .I1(sdpb_inst_15_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(sdpb_inst_16_dout[10]),
  .I1(sdpb_inst_17_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(sdpb_inst_18_dout[10]),
  .I1(sdpb_inst_19_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(sdpb_inst_20_dout[10]),
  .I1(sdpb_inst_21_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(sdpb_inst_22_dout[10]),
  .I1(sdpb_inst_23_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(sdpb_inst_24_dout[10]),
  .I1(sdpb_inst_25_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(sdpb_inst_26_dout[10]),
  .I1(sdpb_inst_27_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(sdpb_inst_28_dout[10]),
  .I1(sdpb_inst_29_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(sdpb_inst_30_dout[10]),
  .I1(sdpb_inst_31_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(sdpb_inst_32_dout[10]),
  .I1(sdpb_inst_33_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(sdpb_inst_34_dout[10]),
  .I1(sdpb_inst_35_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(sdpb_inst_36_dout[10]),
  .I1(sdpb_inst_37_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(sdpb_inst_38_dout[10]),
  .I1(sdpb_inst_39_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(sdpb_inst_40_dout[10]),
  .I1(sdpb_inst_41_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(sdpb_inst_42_dout[10]),
  .I1(sdpb_inst_43_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(sdpb_inst_44_dout[10]),
  .I1(sdpb_inst_45_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(sdpb_inst_46_dout[10]),
  .I1(sdpb_inst_47_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(sdpb_inst_48_dout[10]),
  .I1(sdpb_inst_49_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(sdpb_inst_50_dout[10]),
  .I1(sdpb_inst_51_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(sdpb_inst_52_dout[10]),
  .I1(sdpb_inst_53_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(sdpb_inst_54_dout[10]),
  .I1(sdpb_inst_55_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(sdpb_inst_56_dout[10]),
  .I1(sdpb_inst_57_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(sdpb_inst_58_dout[10]),
  .I1(sdpb_inst_59_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(sdpb_inst_60_dout[10]),
  .I1(sdpb_inst_61_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(sdpb_inst_62_dout[10]),
  .I1(sdpb_inst_63_dout[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(dff_q_4)
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(dff_q_4)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(mux_o_634),
  .I1(mux_o_635),
  .S0(dff_q_4)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(mux_o_636),
  .I1(mux_o_637),
  .S0(dff_q_4)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(dff_q_4)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(mux_o_640),
  .I1(mux_o_641),
  .S0(dff_q_4)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(dff_q_4)
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(mux_o_644),
  .I1(mux_o_645),
  .S0(dff_q_4)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_646),
  .I1(mux_o_647),
  .S0(dff_q_4)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_648),
  .I1(mux_o_649),
  .S0(dff_q_4)
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(mux_o_650),
  .I1(mux_o_651),
  .S0(dff_q_4)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(mux_o_652),
  .I1(mux_o_653),
  .S0(dff_q_4)
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(mux_o_654),
  .I1(mux_o_655),
  .S0(dff_q_4)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(mux_o_656),
  .I1(mux_o_657),
  .S0(dff_q_4)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(mux_o_658),
  .I1(mux_o_659),
  .S0(dff_q_4)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(mux_o_660),
  .I1(mux_o_661),
  .S0(dff_q_4)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(mux_o_662),
  .I1(mux_o_663),
  .S0(dff_q_3)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(mux_o_664),
  .I1(mux_o_665),
  .S0(dff_q_3)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(mux_o_666),
  .I1(mux_o_667),
  .S0(dff_q_3)
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(mux_o_668),
  .I1(mux_o_669),
  .S0(dff_q_3)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(mux_o_670),
  .I1(mux_o_671),
  .S0(dff_q_3)
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(mux_o_672),
  .I1(mux_o_673),
  .S0(dff_q_3)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(mux_o_674),
  .I1(mux_o_675),
  .S0(dff_q_3)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(mux_o_676),
  .I1(mux_o_677),
  .S0(dff_q_3)
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(mux_o_678),
  .I1(mux_o_679),
  .S0(dff_q_2)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(mux_o_680),
  .I1(mux_o_681),
  .S0(dff_q_2)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(mux_o_682),
  .I1(mux_o_683),
  .S0(dff_q_2)
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(dff_q_2)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(mux_o_686),
  .I1(mux_o_687),
  .S0(dff_q_1)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(mux_o_688),
  .I1(mux_o_689),
  .S0(dff_q_1)
);
MUX2 mux_inst_692 (
  .O(dout[10]),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(dff_q_0)
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(sdpb_inst_0_dout[11]),
  .I1(sdpb_inst_1_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(sdpb_inst_2_dout[11]),
  .I1(sdpb_inst_3_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(sdpb_inst_4_dout[11]),
  .I1(sdpb_inst_5_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(sdpb_inst_6_dout[11]),
  .I1(sdpb_inst_7_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(sdpb_inst_8_dout[11]),
  .I1(sdpb_inst_9_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(sdpb_inst_10_dout[11]),
  .I1(sdpb_inst_11_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(sdpb_inst_12_dout[11]),
  .I1(sdpb_inst_13_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(sdpb_inst_14_dout[11]),
  .I1(sdpb_inst_15_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(sdpb_inst_16_dout[11]),
  .I1(sdpb_inst_17_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(sdpb_inst_18_dout[11]),
  .I1(sdpb_inst_19_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(sdpb_inst_20_dout[11]),
  .I1(sdpb_inst_21_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(sdpb_inst_22_dout[11]),
  .I1(sdpb_inst_23_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(sdpb_inst_24_dout[11]),
  .I1(sdpb_inst_25_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(sdpb_inst_26_dout[11]),
  .I1(sdpb_inst_27_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(sdpb_inst_28_dout[11]),
  .I1(sdpb_inst_29_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(sdpb_inst_30_dout[11]),
  .I1(sdpb_inst_31_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(sdpb_inst_32_dout[11]),
  .I1(sdpb_inst_33_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(sdpb_inst_34_dout[11]),
  .I1(sdpb_inst_35_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(sdpb_inst_36_dout[11]),
  .I1(sdpb_inst_37_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(sdpb_inst_38_dout[11]),
  .I1(sdpb_inst_39_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(sdpb_inst_40_dout[11]),
  .I1(sdpb_inst_41_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(sdpb_inst_42_dout[11]),
  .I1(sdpb_inst_43_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(sdpb_inst_44_dout[11]),
  .I1(sdpb_inst_45_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(sdpb_inst_46_dout[11]),
  .I1(sdpb_inst_47_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(sdpb_inst_48_dout[11]),
  .I1(sdpb_inst_49_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(sdpb_inst_50_dout[11]),
  .I1(sdpb_inst_51_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(sdpb_inst_52_dout[11]),
  .I1(sdpb_inst_53_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(sdpb_inst_54_dout[11]),
  .I1(sdpb_inst_55_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(sdpb_inst_56_dout[11]),
  .I1(sdpb_inst_57_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(sdpb_inst_58_dout[11]),
  .I1(sdpb_inst_59_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(sdpb_inst_60_dout[11]),
  .I1(sdpb_inst_61_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(sdpb_inst_62_dout[11]),
  .I1(sdpb_inst_63_dout[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(mux_o_693),
  .I1(mux_o_694),
  .S0(dff_q_4)
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(mux_o_695),
  .I1(mux_o_696),
  .S0(dff_q_4)
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(mux_o_697),
  .I1(mux_o_698),
  .S0(dff_q_4)
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(mux_o_699),
  .I1(mux_o_700),
  .S0(dff_q_4)
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_701),
  .I1(mux_o_702),
  .S0(dff_q_4)
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_703),
  .I1(mux_o_704),
  .S0(dff_q_4)
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(dff_q_4)
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_707),
  .I1(mux_o_708),
  .S0(dff_q_4)
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_709),
  .I1(mux_o_710),
  .S0(dff_q_4)
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_711),
  .I1(mux_o_712),
  .S0(dff_q_4)
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(dff_q_4)
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_4)
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_4)
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(dff_q_4)
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(dff_q_4)
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(dff_q_4)
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_725),
  .I1(mux_o_726),
  .S0(dff_q_3)
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_727),
  .I1(mux_o_728),
  .S0(dff_q_3)
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(dff_q_3)
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(dff_q_3)
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(dff_q_3)
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(dff_q_3)
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(dff_q_3)
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(dff_q_3)
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(dff_q_2)
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(mux_o_743),
  .I1(mux_o_744),
  .S0(dff_q_2)
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(mux_o_745),
  .I1(mux_o_746),
  .S0(dff_q_2)
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(mux_o_747),
  .I1(mux_o_748),
  .S0(dff_q_2)
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(mux_o_749),
  .I1(mux_o_750),
  .S0(dff_q_1)
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(mux_o_751),
  .I1(mux_o_752),
  .S0(dff_q_1)
);
MUX2 mux_inst_755 (
  .O(dout[11]),
  .I0(mux_o_753),
  .I1(mux_o_754),
  .S0(dff_q_0)
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(sdpb_inst_0_dout[12]),
  .I1(sdpb_inst_1_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(sdpb_inst_2_dout[12]),
  .I1(sdpb_inst_3_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(sdpb_inst_4_dout[12]),
  .I1(sdpb_inst_5_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(sdpb_inst_6_dout[12]),
  .I1(sdpb_inst_7_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(sdpb_inst_8_dout[12]),
  .I1(sdpb_inst_9_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(sdpb_inst_10_dout[12]),
  .I1(sdpb_inst_11_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(sdpb_inst_12_dout[12]),
  .I1(sdpb_inst_13_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(sdpb_inst_14_dout[12]),
  .I1(sdpb_inst_15_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(sdpb_inst_16_dout[12]),
  .I1(sdpb_inst_17_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(sdpb_inst_18_dout[12]),
  .I1(sdpb_inst_19_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(sdpb_inst_20_dout[12]),
  .I1(sdpb_inst_21_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(sdpb_inst_22_dout[12]),
  .I1(sdpb_inst_23_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(sdpb_inst_24_dout[12]),
  .I1(sdpb_inst_25_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(sdpb_inst_26_dout[12]),
  .I1(sdpb_inst_27_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(sdpb_inst_28_dout[12]),
  .I1(sdpb_inst_29_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(sdpb_inst_30_dout[12]),
  .I1(sdpb_inst_31_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(sdpb_inst_32_dout[12]),
  .I1(sdpb_inst_33_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(sdpb_inst_34_dout[12]),
  .I1(sdpb_inst_35_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(sdpb_inst_36_dout[12]),
  .I1(sdpb_inst_37_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(sdpb_inst_38_dout[12]),
  .I1(sdpb_inst_39_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(sdpb_inst_40_dout[12]),
  .I1(sdpb_inst_41_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(sdpb_inst_42_dout[12]),
  .I1(sdpb_inst_43_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(sdpb_inst_44_dout[12]),
  .I1(sdpb_inst_45_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(sdpb_inst_46_dout[12]),
  .I1(sdpb_inst_47_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(sdpb_inst_48_dout[12]),
  .I1(sdpb_inst_49_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(sdpb_inst_50_dout[12]),
  .I1(sdpb_inst_51_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(sdpb_inst_52_dout[12]),
  .I1(sdpb_inst_53_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(sdpb_inst_54_dout[12]),
  .I1(sdpb_inst_55_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(sdpb_inst_56_dout[12]),
  .I1(sdpb_inst_57_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(sdpb_inst_58_dout[12]),
  .I1(sdpb_inst_59_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(sdpb_inst_60_dout[12]),
  .I1(sdpb_inst_61_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(sdpb_inst_62_dout[12]),
  .I1(sdpb_inst_63_dout[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(mux_o_756),
  .I1(mux_o_757),
  .S0(dff_q_4)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(mux_o_758),
  .I1(mux_o_759),
  .S0(dff_q_4)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(mux_o_760),
  .I1(mux_o_761),
  .S0(dff_q_4)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(dff_q_4)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(dff_q_4)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(dff_q_4)
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(dff_q_4)
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(dff_q_4)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(dff_q_4)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(mux_o_774),
  .I1(mux_o_775),
  .S0(dff_q_4)
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(mux_o_776),
  .I1(mux_o_777),
  .S0(dff_q_4)
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(mux_o_778),
  .I1(mux_o_779),
  .S0(dff_q_4)
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(mux_o_780),
  .I1(mux_o_781),
  .S0(dff_q_4)
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(mux_o_782),
  .I1(mux_o_783),
  .S0(dff_q_4)
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(mux_o_784),
  .I1(mux_o_785),
  .S0(dff_q_4)
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(mux_o_786),
  .I1(mux_o_787),
  .S0(dff_q_4)
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(mux_o_788),
  .I1(mux_o_789),
  .S0(dff_q_3)
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(mux_o_790),
  .I1(mux_o_791),
  .S0(dff_q_3)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(dff_q_3)
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(mux_o_794),
  .I1(mux_o_795),
  .S0(dff_q_3)
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(mux_o_796),
  .I1(mux_o_797),
  .S0(dff_q_3)
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(mux_o_798),
  .I1(mux_o_799),
  .S0(dff_q_3)
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(mux_o_800),
  .I1(mux_o_801),
  .S0(dff_q_3)
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(mux_o_802),
  .I1(mux_o_803),
  .S0(dff_q_3)
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(mux_o_804),
  .I1(mux_o_805),
  .S0(dff_q_2)
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(dff_q_2)
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(dff_q_2)
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(dff_q_2)
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(dff_q_1)
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(dff_q_1)
);
MUX2 mux_inst_818 (
  .O(dout[12]),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(dff_q_0)
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(sdpb_inst_0_dout[13]),
  .I1(sdpb_inst_1_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(sdpb_inst_2_dout[13]),
  .I1(sdpb_inst_3_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(sdpb_inst_4_dout[13]),
  .I1(sdpb_inst_5_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(sdpb_inst_6_dout[13]),
  .I1(sdpb_inst_7_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(sdpb_inst_8_dout[13]),
  .I1(sdpb_inst_9_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(sdpb_inst_10_dout[13]),
  .I1(sdpb_inst_11_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(sdpb_inst_12_dout[13]),
  .I1(sdpb_inst_13_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(sdpb_inst_14_dout[13]),
  .I1(sdpb_inst_15_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(sdpb_inst_16_dout[13]),
  .I1(sdpb_inst_17_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(sdpb_inst_18_dout[13]),
  .I1(sdpb_inst_19_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(sdpb_inst_20_dout[13]),
  .I1(sdpb_inst_21_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(sdpb_inst_22_dout[13]),
  .I1(sdpb_inst_23_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(sdpb_inst_24_dout[13]),
  .I1(sdpb_inst_25_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(sdpb_inst_26_dout[13]),
  .I1(sdpb_inst_27_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(sdpb_inst_28_dout[13]),
  .I1(sdpb_inst_29_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(sdpb_inst_30_dout[13]),
  .I1(sdpb_inst_31_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(sdpb_inst_32_dout[13]),
  .I1(sdpb_inst_33_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(sdpb_inst_34_dout[13]),
  .I1(sdpb_inst_35_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(sdpb_inst_36_dout[13]),
  .I1(sdpb_inst_37_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(sdpb_inst_38_dout[13]),
  .I1(sdpb_inst_39_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(sdpb_inst_40_dout[13]),
  .I1(sdpb_inst_41_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(sdpb_inst_42_dout[13]),
  .I1(sdpb_inst_43_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(sdpb_inst_44_dout[13]),
  .I1(sdpb_inst_45_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(sdpb_inst_46_dout[13]),
  .I1(sdpb_inst_47_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(sdpb_inst_48_dout[13]),
  .I1(sdpb_inst_49_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(sdpb_inst_50_dout[13]),
  .I1(sdpb_inst_51_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(sdpb_inst_52_dout[13]),
  .I1(sdpb_inst_53_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(sdpb_inst_54_dout[13]),
  .I1(sdpb_inst_55_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(sdpb_inst_56_dout[13]),
  .I1(sdpb_inst_57_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(sdpb_inst_58_dout[13]),
  .I1(sdpb_inst_59_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(sdpb_inst_60_dout[13]),
  .I1(sdpb_inst_61_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(sdpb_inst_62_dout[13]),
  .I1(sdpb_inst_63_dout[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(mux_o_819),
  .I1(mux_o_820),
  .S0(dff_q_4)
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(mux_o_821),
  .I1(mux_o_822),
  .S0(dff_q_4)
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_823),
  .I1(mux_o_824),
  .S0(dff_q_4)
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(mux_o_825),
  .I1(mux_o_826),
  .S0(dff_q_4)
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(mux_o_827),
  .I1(mux_o_828),
  .S0(dff_q_4)
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(mux_o_829),
  .I1(mux_o_830),
  .S0(dff_q_4)
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(mux_o_831),
  .I1(mux_o_832),
  .S0(dff_q_4)
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(mux_o_833),
  .I1(mux_o_834),
  .S0(dff_q_4)
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(mux_o_835),
  .I1(mux_o_836),
  .S0(dff_q_4)
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(mux_o_837),
  .I1(mux_o_838),
  .S0(dff_q_4)
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(mux_o_839),
  .I1(mux_o_840),
  .S0(dff_q_4)
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(mux_o_841),
  .I1(mux_o_842),
  .S0(dff_q_4)
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_843),
  .I1(mux_o_844),
  .S0(dff_q_4)
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_845),
  .I1(mux_o_846),
  .S0(dff_q_4)
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_847),
  .I1(mux_o_848),
  .S0(dff_q_4)
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_849),
  .I1(mux_o_850),
  .S0(dff_q_4)
);
MUX2 mux_inst_867 (
  .O(mux_o_867),
  .I0(mux_o_851),
  .I1(mux_o_852),
  .S0(dff_q_3)
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(mux_o_853),
  .I1(mux_o_854),
  .S0(dff_q_3)
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(mux_o_855),
  .I1(mux_o_856),
  .S0(dff_q_3)
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(mux_o_857),
  .I1(mux_o_858),
  .S0(dff_q_3)
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(mux_o_859),
  .I1(mux_o_860),
  .S0(dff_q_3)
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(mux_o_861),
  .I1(mux_o_862),
  .S0(dff_q_3)
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(mux_o_863),
  .I1(mux_o_864),
  .S0(dff_q_3)
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(mux_o_865),
  .I1(mux_o_866),
  .S0(dff_q_3)
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(mux_o_867),
  .I1(mux_o_868),
  .S0(dff_q_2)
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(mux_o_869),
  .I1(mux_o_870),
  .S0(dff_q_2)
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(mux_o_871),
  .I1(mux_o_872),
  .S0(dff_q_2)
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(mux_o_873),
  .I1(mux_o_874),
  .S0(dff_q_2)
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(mux_o_875),
  .I1(mux_o_876),
  .S0(dff_q_1)
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(mux_o_877),
  .I1(mux_o_878),
  .S0(dff_q_1)
);
MUX2 mux_inst_881 (
  .O(dout[13]),
  .I0(mux_o_879),
  .I1(mux_o_880),
  .S0(dff_q_0)
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(sdpb_inst_0_dout[14]),
  .I1(sdpb_inst_1_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(sdpb_inst_2_dout[14]),
  .I1(sdpb_inst_3_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(sdpb_inst_4_dout[14]),
  .I1(sdpb_inst_5_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(sdpb_inst_6_dout[14]),
  .I1(sdpb_inst_7_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(sdpb_inst_8_dout[14]),
  .I1(sdpb_inst_9_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(sdpb_inst_10_dout[14]),
  .I1(sdpb_inst_11_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_888 (
  .O(mux_o_888),
  .I0(sdpb_inst_12_dout[14]),
  .I1(sdpb_inst_13_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(sdpb_inst_14_dout[14]),
  .I1(sdpb_inst_15_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(sdpb_inst_16_dout[14]),
  .I1(sdpb_inst_17_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(sdpb_inst_18_dout[14]),
  .I1(sdpb_inst_19_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(sdpb_inst_20_dout[14]),
  .I1(sdpb_inst_21_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(sdpb_inst_22_dout[14]),
  .I1(sdpb_inst_23_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(sdpb_inst_24_dout[14]),
  .I1(sdpb_inst_25_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(sdpb_inst_26_dout[14]),
  .I1(sdpb_inst_27_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(sdpb_inst_28_dout[14]),
  .I1(sdpb_inst_29_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(sdpb_inst_30_dout[14]),
  .I1(sdpb_inst_31_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_898 (
  .O(mux_o_898),
  .I0(sdpb_inst_32_dout[14]),
  .I1(sdpb_inst_33_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(sdpb_inst_34_dout[14]),
  .I1(sdpb_inst_35_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(sdpb_inst_36_dout[14]),
  .I1(sdpb_inst_37_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(sdpb_inst_38_dout[14]),
  .I1(sdpb_inst_39_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(sdpb_inst_40_dout[14]),
  .I1(sdpb_inst_41_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(sdpb_inst_42_dout[14]),
  .I1(sdpb_inst_43_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(sdpb_inst_44_dout[14]),
  .I1(sdpb_inst_45_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(sdpb_inst_46_dout[14]),
  .I1(sdpb_inst_47_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(sdpb_inst_48_dout[14]),
  .I1(sdpb_inst_49_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(sdpb_inst_50_dout[14]),
  .I1(sdpb_inst_51_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(sdpb_inst_52_dout[14]),
  .I1(sdpb_inst_53_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(sdpb_inst_54_dout[14]),
  .I1(sdpb_inst_55_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(sdpb_inst_56_dout[14]),
  .I1(sdpb_inst_57_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(sdpb_inst_58_dout[14]),
  .I1(sdpb_inst_59_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(sdpb_inst_60_dout[14]),
  .I1(sdpb_inst_61_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(sdpb_inst_62_dout[14]),
  .I1(sdpb_inst_63_dout[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(dff_q_4)
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(dff_q_4)
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(dff_q_4)
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(mux_o_888),
  .I1(mux_o_889),
  .S0(dff_q_4)
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(mux_o_890),
  .I1(mux_o_891),
  .S0(dff_q_4)
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(mux_o_892),
  .I1(mux_o_893),
  .S0(dff_q_4)
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(mux_o_894),
  .I1(mux_o_895),
  .S0(dff_q_4)
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(mux_o_896),
  .I1(mux_o_897),
  .S0(dff_q_4)
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(mux_o_898),
  .I1(mux_o_899),
  .S0(dff_q_4)
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(mux_o_900),
  .I1(mux_o_901),
  .S0(dff_q_4)
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(mux_o_902),
  .I1(mux_o_903),
  .S0(dff_q_4)
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(mux_o_904),
  .I1(mux_o_905),
  .S0(dff_q_4)
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(mux_o_906),
  .I1(mux_o_907),
  .S0(dff_q_4)
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(mux_o_908),
  .I1(mux_o_909),
  .S0(dff_q_4)
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(mux_o_910),
  .I1(mux_o_911),
  .S0(dff_q_4)
);
MUX2 mux_inst_929 (
  .O(mux_o_929),
  .I0(mux_o_912),
  .I1(mux_o_913),
  .S0(dff_q_4)
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(mux_o_914),
  .I1(mux_o_915),
  .S0(dff_q_3)
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(mux_o_916),
  .I1(mux_o_917),
  .S0(dff_q_3)
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(mux_o_918),
  .I1(mux_o_919),
  .S0(dff_q_3)
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(mux_o_920),
  .I1(mux_o_921),
  .S0(dff_q_3)
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(mux_o_922),
  .I1(mux_o_923),
  .S0(dff_q_3)
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(mux_o_924),
  .I1(mux_o_925),
  .S0(dff_q_3)
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(mux_o_926),
  .I1(mux_o_927),
  .S0(dff_q_3)
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(mux_o_928),
  .I1(mux_o_929),
  .S0(dff_q_3)
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(dff_q_2)
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(dff_q_2)
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(mux_o_934),
  .I1(mux_o_935),
  .S0(dff_q_2)
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(mux_o_936),
  .I1(mux_o_937),
  .S0(dff_q_2)
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(mux_o_938),
  .I1(mux_o_939),
  .S0(dff_q_1)
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(mux_o_940),
  .I1(mux_o_941),
  .S0(dff_q_1)
);
MUX2 mux_inst_944 (
  .O(dout[14]),
  .I0(mux_o_942),
  .I1(mux_o_943),
  .S0(dff_q_0)
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(sdpb_inst_0_dout[15]),
  .I1(sdpb_inst_1_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(sdpb_inst_2_dout[15]),
  .I1(sdpb_inst_3_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(sdpb_inst_4_dout[15]),
  .I1(sdpb_inst_5_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(sdpb_inst_6_dout[15]),
  .I1(sdpb_inst_7_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(sdpb_inst_8_dout[15]),
  .I1(sdpb_inst_9_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(sdpb_inst_10_dout[15]),
  .I1(sdpb_inst_11_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(sdpb_inst_12_dout[15]),
  .I1(sdpb_inst_13_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(sdpb_inst_14_dout[15]),
  .I1(sdpb_inst_15_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(sdpb_inst_16_dout[15]),
  .I1(sdpb_inst_17_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(sdpb_inst_18_dout[15]),
  .I1(sdpb_inst_19_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(sdpb_inst_20_dout[15]),
  .I1(sdpb_inst_21_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(sdpb_inst_22_dout[15]),
  .I1(sdpb_inst_23_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(sdpb_inst_24_dout[15]),
  .I1(sdpb_inst_25_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(sdpb_inst_26_dout[15]),
  .I1(sdpb_inst_27_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(sdpb_inst_28_dout[15]),
  .I1(sdpb_inst_29_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_960 (
  .O(mux_o_960),
  .I0(sdpb_inst_30_dout[15]),
  .I1(sdpb_inst_31_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(sdpb_inst_32_dout[15]),
  .I1(sdpb_inst_33_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(sdpb_inst_34_dout[15]),
  .I1(sdpb_inst_35_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(sdpb_inst_36_dout[15]),
  .I1(sdpb_inst_37_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(sdpb_inst_38_dout[15]),
  .I1(sdpb_inst_39_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(sdpb_inst_40_dout[15]),
  .I1(sdpb_inst_41_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(sdpb_inst_42_dout[15]),
  .I1(sdpb_inst_43_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(sdpb_inst_44_dout[15]),
  .I1(sdpb_inst_45_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(sdpb_inst_46_dout[15]),
  .I1(sdpb_inst_47_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(sdpb_inst_48_dout[15]),
  .I1(sdpb_inst_49_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(sdpb_inst_50_dout[15]),
  .I1(sdpb_inst_51_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(sdpb_inst_52_dout[15]),
  .I1(sdpb_inst_53_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(sdpb_inst_54_dout[15]),
  .I1(sdpb_inst_55_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(sdpb_inst_56_dout[15]),
  .I1(sdpb_inst_57_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(sdpb_inst_58_dout[15]),
  .I1(sdpb_inst_59_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(sdpb_inst_60_dout[15]),
  .I1(sdpb_inst_61_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(sdpb_inst_62_dout[15]),
  .I1(sdpb_inst_63_dout[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(mux_o_945),
  .I1(mux_o_946),
  .S0(dff_q_4)
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(mux_o_947),
  .I1(mux_o_948),
  .S0(dff_q_4)
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(mux_o_949),
  .I1(mux_o_950),
  .S0(dff_q_4)
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(mux_o_951),
  .I1(mux_o_952),
  .S0(dff_q_4)
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(mux_o_953),
  .I1(mux_o_954),
  .S0(dff_q_4)
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(mux_o_955),
  .I1(mux_o_956),
  .S0(dff_q_4)
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(mux_o_957),
  .I1(mux_o_958),
  .S0(dff_q_4)
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(mux_o_959),
  .I1(mux_o_960),
  .S0(dff_q_4)
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(dff_q_4)
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(dff_q_4)
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(dff_q_4)
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(mux_o_967),
  .I1(mux_o_968),
  .S0(dff_q_4)
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(mux_o_969),
  .I1(mux_o_970),
  .S0(dff_q_4)
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(mux_o_971),
  .I1(mux_o_972),
  .S0(dff_q_4)
);
MUX2 mux_inst_991 (
  .O(mux_o_991),
  .I0(mux_o_973),
  .I1(mux_o_974),
  .S0(dff_q_4)
);
MUX2 mux_inst_992 (
  .O(mux_o_992),
  .I0(mux_o_975),
  .I1(mux_o_976),
  .S0(dff_q_4)
);
MUX2 mux_inst_993 (
  .O(mux_o_993),
  .I0(mux_o_977),
  .I1(mux_o_978),
  .S0(dff_q_3)
);
MUX2 mux_inst_994 (
  .O(mux_o_994),
  .I0(mux_o_979),
  .I1(mux_o_980),
  .S0(dff_q_3)
);
MUX2 mux_inst_995 (
  .O(mux_o_995),
  .I0(mux_o_981),
  .I1(mux_o_982),
  .S0(dff_q_3)
);
MUX2 mux_inst_996 (
  .O(mux_o_996),
  .I0(mux_o_983),
  .I1(mux_o_984),
  .S0(dff_q_3)
);
MUX2 mux_inst_997 (
  .O(mux_o_997),
  .I0(mux_o_985),
  .I1(mux_o_986),
  .S0(dff_q_3)
);
MUX2 mux_inst_998 (
  .O(mux_o_998),
  .I0(mux_o_987),
  .I1(mux_o_988),
  .S0(dff_q_3)
);
MUX2 mux_inst_999 (
  .O(mux_o_999),
  .I0(mux_o_989),
  .I1(mux_o_990),
  .S0(dff_q_3)
);
MUX2 mux_inst_1000 (
  .O(mux_o_1000),
  .I0(mux_o_991),
  .I1(mux_o_992),
  .S0(dff_q_3)
);
MUX2 mux_inst_1001 (
  .O(mux_o_1001),
  .I0(mux_o_993),
  .I1(mux_o_994),
  .S0(dff_q_2)
);
MUX2 mux_inst_1002 (
  .O(mux_o_1002),
  .I0(mux_o_995),
  .I1(mux_o_996),
  .S0(dff_q_2)
);
MUX2 mux_inst_1003 (
  .O(mux_o_1003),
  .I0(mux_o_997),
  .I1(mux_o_998),
  .S0(dff_q_2)
);
MUX2 mux_inst_1004 (
  .O(mux_o_1004),
  .I0(mux_o_999),
  .I1(mux_o_1000),
  .S0(dff_q_2)
);
MUX2 mux_inst_1005 (
  .O(mux_o_1005),
  .I0(mux_o_1001),
  .I1(mux_o_1002),
  .S0(dff_q_1)
);
MUX2 mux_inst_1006 (
  .O(mux_o_1006),
  .I0(mux_o_1003),
  .I1(mux_o_1004),
  .S0(dff_q_1)
);
MUX2 mux_inst_1007 (
  .O(dout[15]),
  .I0(mux_o_1005),
  .I1(mux_o_1006),
  .S0(dff_q_0)
);
MUX2 mux_inst_1008 (
  .O(mux_o_1008),
  .I0(sdpb_inst_64_dout[16]),
  .I1(sdpb_inst_65_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1009 (
  .O(mux_o_1009),
  .I0(sdpb_inst_66_dout[16]),
  .I1(sdpb_inst_67_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1010 (
  .O(mux_o_1010),
  .I0(sdpb_inst_68_dout[16]),
  .I1(sdpb_inst_69_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1011 (
  .O(mux_o_1011),
  .I0(sdpb_inst_70_dout[16]),
  .I1(sdpb_inst_71_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1012 (
  .O(mux_o_1012),
  .I0(sdpb_inst_72_dout[16]),
  .I1(sdpb_inst_73_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1013 (
  .O(mux_o_1013),
  .I0(sdpb_inst_74_dout[16]),
  .I1(sdpb_inst_75_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1014 (
  .O(mux_o_1014),
  .I0(sdpb_inst_76_dout[16]),
  .I1(sdpb_inst_77_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1015 (
  .O(mux_o_1015),
  .I0(sdpb_inst_78_dout[16]),
  .I1(sdpb_inst_79_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1016 (
  .O(mux_o_1016),
  .I0(sdpb_inst_80_dout[16]),
  .I1(sdpb_inst_81_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1017 (
  .O(mux_o_1017),
  .I0(sdpb_inst_82_dout[16]),
  .I1(sdpb_inst_83_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1018 (
  .O(mux_o_1018),
  .I0(sdpb_inst_84_dout[16]),
  .I1(sdpb_inst_85_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1019 (
  .O(mux_o_1019),
  .I0(sdpb_inst_86_dout[16]),
  .I1(sdpb_inst_87_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1020 (
  .O(mux_o_1020),
  .I0(sdpb_inst_88_dout[16]),
  .I1(sdpb_inst_89_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1021 (
  .O(mux_o_1021),
  .I0(sdpb_inst_90_dout[16]),
  .I1(sdpb_inst_91_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1022 (
  .O(mux_o_1022),
  .I0(sdpb_inst_92_dout[16]),
  .I1(sdpb_inst_93_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1023 (
  .O(mux_o_1023),
  .I0(sdpb_inst_94_dout[16]),
  .I1(sdpb_inst_95_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1024 (
  .O(mux_o_1024),
  .I0(sdpb_inst_96_dout[16]),
  .I1(sdpb_inst_97_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1025 (
  .O(mux_o_1025),
  .I0(sdpb_inst_98_dout[16]),
  .I1(sdpb_inst_99_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1026 (
  .O(mux_o_1026),
  .I0(sdpb_inst_100_dout[16]),
  .I1(sdpb_inst_101_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1027 (
  .O(mux_o_1027),
  .I0(sdpb_inst_102_dout[16]),
  .I1(sdpb_inst_103_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1028 (
  .O(mux_o_1028),
  .I0(sdpb_inst_104_dout[16]),
  .I1(sdpb_inst_105_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1029 (
  .O(mux_o_1029),
  .I0(sdpb_inst_106_dout[16]),
  .I1(sdpb_inst_107_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1030 (
  .O(mux_o_1030),
  .I0(sdpb_inst_108_dout[16]),
  .I1(sdpb_inst_109_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1031 (
  .O(mux_o_1031),
  .I0(sdpb_inst_110_dout[16]),
  .I1(sdpb_inst_111_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1032 (
  .O(mux_o_1032),
  .I0(sdpb_inst_112_dout[16]),
  .I1(sdpb_inst_113_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1033 (
  .O(mux_o_1033),
  .I0(sdpb_inst_114_dout[16]),
  .I1(sdpb_inst_115_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1034 (
  .O(mux_o_1034),
  .I0(sdpb_inst_116_dout[16]),
  .I1(sdpb_inst_117_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1035 (
  .O(mux_o_1035),
  .I0(sdpb_inst_118_dout[16]),
  .I1(sdpb_inst_119_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1036 (
  .O(mux_o_1036),
  .I0(sdpb_inst_120_dout[16]),
  .I1(sdpb_inst_121_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1037 (
  .O(mux_o_1037),
  .I0(sdpb_inst_122_dout[16]),
  .I1(sdpb_inst_123_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1038 (
  .O(mux_o_1038),
  .I0(sdpb_inst_124_dout[16]),
  .I1(sdpb_inst_125_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1039 (
  .O(mux_o_1039),
  .I0(sdpb_inst_126_dout[16]),
  .I1(sdpb_inst_127_dout[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1040 (
  .O(mux_o_1040),
  .I0(mux_o_1008),
  .I1(mux_o_1009),
  .S0(dff_q_4)
);
MUX2 mux_inst_1041 (
  .O(mux_o_1041),
  .I0(mux_o_1010),
  .I1(mux_o_1011),
  .S0(dff_q_4)
);
MUX2 mux_inst_1042 (
  .O(mux_o_1042),
  .I0(mux_o_1012),
  .I1(mux_o_1013),
  .S0(dff_q_4)
);
MUX2 mux_inst_1043 (
  .O(mux_o_1043),
  .I0(mux_o_1014),
  .I1(mux_o_1015),
  .S0(dff_q_4)
);
MUX2 mux_inst_1044 (
  .O(mux_o_1044),
  .I0(mux_o_1016),
  .I1(mux_o_1017),
  .S0(dff_q_4)
);
MUX2 mux_inst_1045 (
  .O(mux_o_1045),
  .I0(mux_o_1018),
  .I1(mux_o_1019),
  .S0(dff_q_4)
);
MUX2 mux_inst_1046 (
  .O(mux_o_1046),
  .I0(mux_o_1020),
  .I1(mux_o_1021),
  .S0(dff_q_4)
);
MUX2 mux_inst_1047 (
  .O(mux_o_1047),
  .I0(mux_o_1022),
  .I1(mux_o_1023),
  .S0(dff_q_4)
);
MUX2 mux_inst_1048 (
  .O(mux_o_1048),
  .I0(mux_o_1024),
  .I1(mux_o_1025),
  .S0(dff_q_4)
);
MUX2 mux_inst_1049 (
  .O(mux_o_1049),
  .I0(mux_o_1026),
  .I1(mux_o_1027),
  .S0(dff_q_4)
);
MUX2 mux_inst_1050 (
  .O(mux_o_1050),
  .I0(mux_o_1028),
  .I1(mux_o_1029),
  .S0(dff_q_4)
);
MUX2 mux_inst_1051 (
  .O(mux_o_1051),
  .I0(mux_o_1030),
  .I1(mux_o_1031),
  .S0(dff_q_4)
);
MUX2 mux_inst_1052 (
  .O(mux_o_1052),
  .I0(mux_o_1032),
  .I1(mux_o_1033),
  .S0(dff_q_4)
);
MUX2 mux_inst_1053 (
  .O(mux_o_1053),
  .I0(mux_o_1034),
  .I1(mux_o_1035),
  .S0(dff_q_4)
);
MUX2 mux_inst_1054 (
  .O(mux_o_1054),
  .I0(mux_o_1036),
  .I1(mux_o_1037),
  .S0(dff_q_4)
);
MUX2 mux_inst_1055 (
  .O(mux_o_1055),
  .I0(mux_o_1038),
  .I1(mux_o_1039),
  .S0(dff_q_4)
);
MUX2 mux_inst_1056 (
  .O(mux_o_1056),
  .I0(mux_o_1040),
  .I1(mux_o_1041),
  .S0(dff_q_3)
);
MUX2 mux_inst_1057 (
  .O(mux_o_1057),
  .I0(mux_o_1042),
  .I1(mux_o_1043),
  .S0(dff_q_3)
);
MUX2 mux_inst_1058 (
  .O(mux_o_1058),
  .I0(mux_o_1044),
  .I1(mux_o_1045),
  .S0(dff_q_3)
);
MUX2 mux_inst_1059 (
  .O(mux_o_1059),
  .I0(mux_o_1046),
  .I1(mux_o_1047),
  .S0(dff_q_3)
);
MUX2 mux_inst_1060 (
  .O(mux_o_1060),
  .I0(mux_o_1048),
  .I1(mux_o_1049),
  .S0(dff_q_3)
);
MUX2 mux_inst_1061 (
  .O(mux_o_1061),
  .I0(mux_o_1050),
  .I1(mux_o_1051),
  .S0(dff_q_3)
);
MUX2 mux_inst_1062 (
  .O(mux_o_1062),
  .I0(mux_o_1052),
  .I1(mux_o_1053),
  .S0(dff_q_3)
);
MUX2 mux_inst_1063 (
  .O(mux_o_1063),
  .I0(mux_o_1054),
  .I1(mux_o_1055),
  .S0(dff_q_3)
);
MUX2 mux_inst_1064 (
  .O(mux_o_1064),
  .I0(mux_o_1056),
  .I1(mux_o_1057),
  .S0(dff_q_2)
);
MUX2 mux_inst_1065 (
  .O(mux_o_1065),
  .I0(mux_o_1058),
  .I1(mux_o_1059),
  .S0(dff_q_2)
);
MUX2 mux_inst_1066 (
  .O(mux_o_1066),
  .I0(mux_o_1060),
  .I1(mux_o_1061),
  .S0(dff_q_2)
);
MUX2 mux_inst_1067 (
  .O(mux_o_1067),
  .I0(mux_o_1062),
  .I1(mux_o_1063),
  .S0(dff_q_2)
);
MUX2 mux_inst_1068 (
  .O(mux_o_1068),
  .I0(mux_o_1064),
  .I1(mux_o_1065),
  .S0(dff_q_1)
);
MUX2 mux_inst_1069 (
  .O(mux_o_1069),
  .I0(mux_o_1066),
  .I1(mux_o_1067),
  .S0(dff_q_1)
);
MUX2 mux_inst_1070 (
  .O(dout[16]),
  .I0(mux_o_1068),
  .I1(mux_o_1069),
  .S0(dff_q_0)
);
MUX2 mux_inst_1071 (
  .O(mux_o_1071),
  .I0(sdpb_inst_64_dout[17]),
  .I1(sdpb_inst_65_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1072 (
  .O(mux_o_1072),
  .I0(sdpb_inst_66_dout[17]),
  .I1(sdpb_inst_67_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1073 (
  .O(mux_o_1073),
  .I0(sdpb_inst_68_dout[17]),
  .I1(sdpb_inst_69_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1074 (
  .O(mux_o_1074),
  .I0(sdpb_inst_70_dout[17]),
  .I1(sdpb_inst_71_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1075 (
  .O(mux_o_1075),
  .I0(sdpb_inst_72_dout[17]),
  .I1(sdpb_inst_73_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1076 (
  .O(mux_o_1076),
  .I0(sdpb_inst_74_dout[17]),
  .I1(sdpb_inst_75_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1077 (
  .O(mux_o_1077),
  .I0(sdpb_inst_76_dout[17]),
  .I1(sdpb_inst_77_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1078 (
  .O(mux_o_1078),
  .I0(sdpb_inst_78_dout[17]),
  .I1(sdpb_inst_79_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1079 (
  .O(mux_o_1079),
  .I0(sdpb_inst_80_dout[17]),
  .I1(sdpb_inst_81_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1080 (
  .O(mux_o_1080),
  .I0(sdpb_inst_82_dout[17]),
  .I1(sdpb_inst_83_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1081 (
  .O(mux_o_1081),
  .I0(sdpb_inst_84_dout[17]),
  .I1(sdpb_inst_85_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1082 (
  .O(mux_o_1082),
  .I0(sdpb_inst_86_dout[17]),
  .I1(sdpb_inst_87_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1083 (
  .O(mux_o_1083),
  .I0(sdpb_inst_88_dout[17]),
  .I1(sdpb_inst_89_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1084 (
  .O(mux_o_1084),
  .I0(sdpb_inst_90_dout[17]),
  .I1(sdpb_inst_91_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1085 (
  .O(mux_o_1085),
  .I0(sdpb_inst_92_dout[17]),
  .I1(sdpb_inst_93_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1086 (
  .O(mux_o_1086),
  .I0(sdpb_inst_94_dout[17]),
  .I1(sdpb_inst_95_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1087 (
  .O(mux_o_1087),
  .I0(sdpb_inst_96_dout[17]),
  .I1(sdpb_inst_97_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1088 (
  .O(mux_o_1088),
  .I0(sdpb_inst_98_dout[17]),
  .I1(sdpb_inst_99_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1089 (
  .O(mux_o_1089),
  .I0(sdpb_inst_100_dout[17]),
  .I1(sdpb_inst_101_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1090 (
  .O(mux_o_1090),
  .I0(sdpb_inst_102_dout[17]),
  .I1(sdpb_inst_103_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1091 (
  .O(mux_o_1091),
  .I0(sdpb_inst_104_dout[17]),
  .I1(sdpb_inst_105_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1092 (
  .O(mux_o_1092),
  .I0(sdpb_inst_106_dout[17]),
  .I1(sdpb_inst_107_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1093 (
  .O(mux_o_1093),
  .I0(sdpb_inst_108_dout[17]),
  .I1(sdpb_inst_109_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1094 (
  .O(mux_o_1094),
  .I0(sdpb_inst_110_dout[17]),
  .I1(sdpb_inst_111_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1095 (
  .O(mux_o_1095),
  .I0(sdpb_inst_112_dout[17]),
  .I1(sdpb_inst_113_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1096 (
  .O(mux_o_1096),
  .I0(sdpb_inst_114_dout[17]),
  .I1(sdpb_inst_115_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1097 (
  .O(mux_o_1097),
  .I0(sdpb_inst_116_dout[17]),
  .I1(sdpb_inst_117_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1098 (
  .O(mux_o_1098),
  .I0(sdpb_inst_118_dout[17]),
  .I1(sdpb_inst_119_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1099 (
  .O(mux_o_1099),
  .I0(sdpb_inst_120_dout[17]),
  .I1(sdpb_inst_121_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1100 (
  .O(mux_o_1100),
  .I0(sdpb_inst_122_dout[17]),
  .I1(sdpb_inst_123_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1101 (
  .O(mux_o_1101),
  .I0(sdpb_inst_124_dout[17]),
  .I1(sdpb_inst_125_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1102 (
  .O(mux_o_1102),
  .I0(sdpb_inst_126_dout[17]),
  .I1(sdpb_inst_127_dout[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1103 (
  .O(mux_o_1103),
  .I0(mux_o_1071),
  .I1(mux_o_1072),
  .S0(dff_q_4)
);
MUX2 mux_inst_1104 (
  .O(mux_o_1104),
  .I0(mux_o_1073),
  .I1(mux_o_1074),
  .S0(dff_q_4)
);
MUX2 mux_inst_1105 (
  .O(mux_o_1105),
  .I0(mux_o_1075),
  .I1(mux_o_1076),
  .S0(dff_q_4)
);
MUX2 mux_inst_1106 (
  .O(mux_o_1106),
  .I0(mux_o_1077),
  .I1(mux_o_1078),
  .S0(dff_q_4)
);
MUX2 mux_inst_1107 (
  .O(mux_o_1107),
  .I0(mux_o_1079),
  .I1(mux_o_1080),
  .S0(dff_q_4)
);
MUX2 mux_inst_1108 (
  .O(mux_o_1108),
  .I0(mux_o_1081),
  .I1(mux_o_1082),
  .S0(dff_q_4)
);
MUX2 mux_inst_1109 (
  .O(mux_o_1109),
  .I0(mux_o_1083),
  .I1(mux_o_1084),
  .S0(dff_q_4)
);
MUX2 mux_inst_1110 (
  .O(mux_o_1110),
  .I0(mux_o_1085),
  .I1(mux_o_1086),
  .S0(dff_q_4)
);
MUX2 mux_inst_1111 (
  .O(mux_o_1111),
  .I0(mux_o_1087),
  .I1(mux_o_1088),
  .S0(dff_q_4)
);
MUX2 mux_inst_1112 (
  .O(mux_o_1112),
  .I0(mux_o_1089),
  .I1(mux_o_1090),
  .S0(dff_q_4)
);
MUX2 mux_inst_1113 (
  .O(mux_o_1113),
  .I0(mux_o_1091),
  .I1(mux_o_1092),
  .S0(dff_q_4)
);
MUX2 mux_inst_1114 (
  .O(mux_o_1114),
  .I0(mux_o_1093),
  .I1(mux_o_1094),
  .S0(dff_q_4)
);
MUX2 mux_inst_1115 (
  .O(mux_o_1115),
  .I0(mux_o_1095),
  .I1(mux_o_1096),
  .S0(dff_q_4)
);
MUX2 mux_inst_1116 (
  .O(mux_o_1116),
  .I0(mux_o_1097),
  .I1(mux_o_1098),
  .S0(dff_q_4)
);
MUX2 mux_inst_1117 (
  .O(mux_o_1117),
  .I0(mux_o_1099),
  .I1(mux_o_1100),
  .S0(dff_q_4)
);
MUX2 mux_inst_1118 (
  .O(mux_o_1118),
  .I0(mux_o_1101),
  .I1(mux_o_1102),
  .S0(dff_q_4)
);
MUX2 mux_inst_1119 (
  .O(mux_o_1119),
  .I0(mux_o_1103),
  .I1(mux_o_1104),
  .S0(dff_q_3)
);
MUX2 mux_inst_1120 (
  .O(mux_o_1120),
  .I0(mux_o_1105),
  .I1(mux_o_1106),
  .S0(dff_q_3)
);
MUX2 mux_inst_1121 (
  .O(mux_o_1121),
  .I0(mux_o_1107),
  .I1(mux_o_1108),
  .S0(dff_q_3)
);
MUX2 mux_inst_1122 (
  .O(mux_o_1122),
  .I0(mux_o_1109),
  .I1(mux_o_1110),
  .S0(dff_q_3)
);
MUX2 mux_inst_1123 (
  .O(mux_o_1123),
  .I0(mux_o_1111),
  .I1(mux_o_1112),
  .S0(dff_q_3)
);
MUX2 mux_inst_1124 (
  .O(mux_o_1124),
  .I0(mux_o_1113),
  .I1(mux_o_1114),
  .S0(dff_q_3)
);
MUX2 mux_inst_1125 (
  .O(mux_o_1125),
  .I0(mux_o_1115),
  .I1(mux_o_1116),
  .S0(dff_q_3)
);
MUX2 mux_inst_1126 (
  .O(mux_o_1126),
  .I0(mux_o_1117),
  .I1(mux_o_1118),
  .S0(dff_q_3)
);
MUX2 mux_inst_1127 (
  .O(mux_o_1127),
  .I0(mux_o_1119),
  .I1(mux_o_1120),
  .S0(dff_q_2)
);
MUX2 mux_inst_1128 (
  .O(mux_o_1128),
  .I0(mux_o_1121),
  .I1(mux_o_1122),
  .S0(dff_q_2)
);
MUX2 mux_inst_1129 (
  .O(mux_o_1129),
  .I0(mux_o_1123),
  .I1(mux_o_1124),
  .S0(dff_q_2)
);
MUX2 mux_inst_1130 (
  .O(mux_o_1130),
  .I0(mux_o_1125),
  .I1(mux_o_1126),
  .S0(dff_q_2)
);
MUX2 mux_inst_1131 (
  .O(mux_o_1131),
  .I0(mux_o_1127),
  .I1(mux_o_1128),
  .S0(dff_q_1)
);
MUX2 mux_inst_1132 (
  .O(mux_o_1132),
  .I0(mux_o_1129),
  .I1(mux_o_1130),
  .S0(dff_q_1)
);
MUX2 mux_inst_1133 (
  .O(dout[17]),
  .I0(mux_o_1131),
  .I1(mux_o_1132),
  .S0(dff_q_0)
);
MUX2 mux_inst_1134 (
  .O(mux_o_1134),
  .I0(sdpb_inst_64_dout[18]),
  .I1(sdpb_inst_65_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1135 (
  .O(mux_o_1135),
  .I0(sdpb_inst_66_dout[18]),
  .I1(sdpb_inst_67_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1136 (
  .O(mux_o_1136),
  .I0(sdpb_inst_68_dout[18]),
  .I1(sdpb_inst_69_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1137 (
  .O(mux_o_1137),
  .I0(sdpb_inst_70_dout[18]),
  .I1(sdpb_inst_71_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1138 (
  .O(mux_o_1138),
  .I0(sdpb_inst_72_dout[18]),
  .I1(sdpb_inst_73_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1139 (
  .O(mux_o_1139),
  .I0(sdpb_inst_74_dout[18]),
  .I1(sdpb_inst_75_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1140 (
  .O(mux_o_1140),
  .I0(sdpb_inst_76_dout[18]),
  .I1(sdpb_inst_77_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1141 (
  .O(mux_o_1141),
  .I0(sdpb_inst_78_dout[18]),
  .I1(sdpb_inst_79_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1142 (
  .O(mux_o_1142),
  .I0(sdpb_inst_80_dout[18]),
  .I1(sdpb_inst_81_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1143 (
  .O(mux_o_1143),
  .I0(sdpb_inst_82_dout[18]),
  .I1(sdpb_inst_83_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1144 (
  .O(mux_o_1144),
  .I0(sdpb_inst_84_dout[18]),
  .I1(sdpb_inst_85_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1145 (
  .O(mux_o_1145),
  .I0(sdpb_inst_86_dout[18]),
  .I1(sdpb_inst_87_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1146 (
  .O(mux_o_1146),
  .I0(sdpb_inst_88_dout[18]),
  .I1(sdpb_inst_89_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1147 (
  .O(mux_o_1147),
  .I0(sdpb_inst_90_dout[18]),
  .I1(sdpb_inst_91_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1148 (
  .O(mux_o_1148),
  .I0(sdpb_inst_92_dout[18]),
  .I1(sdpb_inst_93_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1149 (
  .O(mux_o_1149),
  .I0(sdpb_inst_94_dout[18]),
  .I1(sdpb_inst_95_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1150 (
  .O(mux_o_1150),
  .I0(sdpb_inst_96_dout[18]),
  .I1(sdpb_inst_97_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1151 (
  .O(mux_o_1151),
  .I0(sdpb_inst_98_dout[18]),
  .I1(sdpb_inst_99_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1152 (
  .O(mux_o_1152),
  .I0(sdpb_inst_100_dout[18]),
  .I1(sdpb_inst_101_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1153 (
  .O(mux_o_1153),
  .I0(sdpb_inst_102_dout[18]),
  .I1(sdpb_inst_103_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1154 (
  .O(mux_o_1154),
  .I0(sdpb_inst_104_dout[18]),
  .I1(sdpb_inst_105_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1155 (
  .O(mux_o_1155),
  .I0(sdpb_inst_106_dout[18]),
  .I1(sdpb_inst_107_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1156 (
  .O(mux_o_1156),
  .I0(sdpb_inst_108_dout[18]),
  .I1(sdpb_inst_109_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1157 (
  .O(mux_o_1157),
  .I0(sdpb_inst_110_dout[18]),
  .I1(sdpb_inst_111_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1158 (
  .O(mux_o_1158),
  .I0(sdpb_inst_112_dout[18]),
  .I1(sdpb_inst_113_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1159 (
  .O(mux_o_1159),
  .I0(sdpb_inst_114_dout[18]),
  .I1(sdpb_inst_115_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1160 (
  .O(mux_o_1160),
  .I0(sdpb_inst_116_dout[18]),
  .I1(sdpb_inst_117_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1161 (
  .O(mux_o_1161),
  .I0(sdpb_inst_118_dout[18]),
  .I1(sdpb_inst_119_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1162 (
  .O(mux_o_1162),
  .I0(sdpb_inst_120_dout[18]),
  .I1(sdpb_inst_121_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1163 (
  .O(mux_o_1163),
  .I0(sdpb_inst_122_dout[18]),
  .I1(sdpb_inst_123_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1164 (
  .O(mux_o_1164),
  .I0(sdpb_inst_124_dout[18]),
  .I1(sdpb_inst_125_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1165 (
  .O(mux_o_1165),
  .I0(sdpb_inst_126_dout[18]),
  .I1(sdpb_inst_127_dout[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1166 (
  .O(mux_o_1166),
  .I0(mux_o_1134),
  .I1(mux_o_1135),
  .S0(dff_q_4)
);
MUX2 mux_inst_1167 (
  .O(mux_o_1167),
  .I0(mux_o_1136),
  .I1(mux_o_1137),
  .S0(dff_q_4)
);
MUX2 mux_inst_1168 (
  .O(mux_o_1168),
  .I0(mux_o_1138),
  .I1(mux_o_1139),
  .S0(dff_q_4)
);
MUX2 mux_inst_1169 (
  .O(mux_o_1169),
  .I0(mux_o_1140),
  .I1(mux_o_1141),
  .S0(dff_q_4)
);
MUX2 mux_inst_1170 (
  .O(mux_o_1170),
  .I0(mux_o_1142),
  .I1(mux_o_1143),
  .S0(dff_q_4)
);
MUX2 mux_inst_1171 (
  .O(mux_o_1171),
  .I0(mux_o_1144),
  .I1(mux_o_1145),
  .S0(dff_q_4)
);
MUX2 mux_inst_1172 (
  .O(mux_o_1172),
  .I0(mux_o_1146),
  .I1(mux_o_1147),
  .S0(dff_q_4)
);
MUX2 mux_inst_1173 (
  .O(mux_o_1173),
  .I0(mux_o_1148),
  .I1(mux_o_1149),
  .S0(dff_q_4)
);
MUX2 mux_inst_1174 (
  .O(mux_o_1174),
  .I0(mux_o_1150),
  .I1(mux_o_1151),
  .S0(dff_q_4)
);
MUX2 mux_inst_1175 (
  .O(mux_o_1175),
  .I0(mux_o_1152),
  .I1(mux_o_1153),
  .S0(dff_q_4)
);
MUX2 mux_inst_1176 (
  .O(mux_o_1176),
  .I0(mux_o_1154),
  .I1(mux_o_1155),
  .S0(dff_q_4)
);
MUX2 mux_inst_1177 (
  .O(mux_o_1177),
  .I0(mux_o_1156),
  .I1(mux_o_1157),
  .S0(dff_q_4)
);
MUX2 mux_inst_1178 (
  .O(mux_o_1178),
  .I0(mux_o_1158),
  .I1(mux_o_1159),
  .S0(dff_q_4)
);
MUX2 mux_inst_1179 (
  .O(mux_o_1179),
  .I0(mux_o_1160),
  .I1(mux_o_1161),
  .S0(dff_q_4)
);
MUX2 mux_inst_1180 (
  .O(mux_o_1180),
  .I0(mux_o_1162),
  .I1(mux_o_1163),
  .S0(dff_q_4)
);
MUX2 mux_inst_1181 (
  .O(mux_o_1181),
  .I0(mux_o_1164),
  .I1(mux_o_1165),
  .S0(dff_q_4)
);
MUX2 mux_inst_1182 (
  .O(mux_o_1182),
  .I0(mux_o_1166),
  .I1(mux_o_1167),
  .S0(dff_q_3)
);
MUX2 mux_inst_1183 (
  .O(mux_o_1183),
  .I0(mux_o_1168),
  .I1(mux_o_1169),
  .S0(dff_q_3)
);
MUX2 mux_inst_1184 (
  .O(mux_o_1184),
  .I0(mux_o_1170),
  .I1(mux_o_1171),
  .S0(dff_q_3)
);
MUX2 mux_inst_1185 (
  .O(mux_o_1185),
  .I0(mux_o_1172),
  .I1(mux_o_1173),
  .S0(dff_q_3)
);
MUX2 mux_inst_1186 (
  .O(mux_o_1186),
  .I0(mux_o_1174),
  .I1(mux_o_1175),
  .S0(dff_q_3)
);
MUX2 mux_inst_1187 (
  .O(mux_o_1187),
  .I0(mux_o_1176),
  .I1(mux_o_1177),
  .S0(dff_q_3)
);
MUX2 mux_inst_1188 (
  .O(mux_o_1188),
  .I0(mux_o_1178),
  .I1(mux_o_1179),
  .S0(dff_q_3)
);
MUX2 mux_inst_1189 (
  .O(mux_o_1189),
  .I0(mux_o_1180),
  .I1(mux_o_1181),
  .S0(dff_q_3)
);
MUX2 mux_inst_1190 (
  .O(mux_o_1190),
  .I0(mux_o_1182),
  .I1(mux_o_1183),
  .S0(dff_q_2)
);
MUX2 mux_inst_1191 (
  .O(mux_o_1191),
  .I0(mux_o_1184),
  .I1(mux_o_1185),
  .S0(dff_q_2)
);
MUX2 mux_inst_1192 (
  .O(mux_o_1192),
  .I0(mux_o_1186),
  .I1(mux_o_1187),
  .S0(dff_q_2)
);
MUX2 mux_inst_1193 (
  .O(mux_o_1193),
  .I0(mux_o_1188),
  .I1(mux_o_1189),
  .S0(dff_q_2)
);
MUX2 mux_inst_1194 (
  .O(mux_o_1194),
  .I0(mux_o_1190),
  .I1(mux_o_1191),
  .S0(dff_q_1)
);
MUX2 mux_inst_1195 (
  .O(mux_o_1195),
  .I0(mux_o_1192),
  .I1(mux_o_1193),
  .S0(dff_q_1)
);
MUX2 mux_inst_1196 (
  .O(dout[18]),
  .I0(mux_o_1194),
  .I1(mux_o_1195),
  .S0(dff_q_0)
);
MUX2 mux_inst_1197 (
  .O(mux_o_1197),
  .I0(sdpb_inst_64_dout[19]),
  .I1(sdpb_inst_65_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1198 (
  .O(mux_o_1198),
  .I0(sdpb_inst_66_dout[19]),
  .I1(sdpb_inst_67_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1199 (
  .O(mux_o_1199),
  .I0(sdpb_inst_68_dout[19]),
  .I1(sdpb_inst_69_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1200 (
  .O(mux_o_1200),
  .I0(sdpb_inst_70_dout[19]),
  .I1(sdpb_inst_71_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1201 (
  .O(mux_o_1201),
  .I0(sdpb_inst_72_dout[19]),
  .I1(sdpb_inst_73_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1202 (
  .O(mux_o_1202),
  .I0(sdpb_inst_74_dout[19]),
  .I1(sdpb_inst_75_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1203 (
  .O(mux_o_1203),
  .I0(sdpb_inst_76_dout[19]),
  .I1(sdpb_inst_77_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1204 (
  .O(mux_o_1204),
  .I0(sdpb_inst_78_dout[19]),
  .I1(sdpb_inst_79_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1205 (
  .O(mux_o_1205),
  .I0(sdpb_inst_80_dout[19]),
  .I1(sdpb_inst_81_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1206 (
  .O(mux_o_1206),
  .I0(sdpb_inst_82_dout[19]),
  .I1(sdpb_inst_83_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1207 (
  .O(mux_o_1207),
  .I0(sdpb_inst_84_dout[19]),
  .I1(sdpb_inst_85_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1208 (
  .O(mux_o_1208),
  .I0(sdpb_inst_86_dout[19]),
  .I1(sdpb_inst_87_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1209 (
  .O(mux_o_1209),
  .I0(sdpb_inst_88_dout[19]),
  .I1(sdpb_inst_89_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1210 (
  .O(mux_o_1210),
  .I0(sdpb_inst_90_dout[19]),
  .I1(sdpb_inst_91_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1211 (
  .O(mux_o_1211),
  .I0(sdpb_inst_92_dout[19]),
  .I1(sdpb_inst_93_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1212 (
  .O(mux_o_1212),
  .I0(sdpb_inst_94_dout[19]),
  .I1(sdpb_inst_95_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1213 (
  .O(mux_o_1213),
  .I0(sdpb_inst_96_dout[19]),
  .I1(sdpb_inst_97_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1214 (
  .O(mux_o_1214),
  .I0(sdpb_inst_98_dout[19]),
  .I1(sdpb_inst_99_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1215 (
  .O(mux_o_1215),
  .I0(sdpb_inst_100_dout[19]),
  .I1(sdpb_inst_101_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1216 (
  .O(mux_o_1216),
  .I0(sdpb_inst_102_dout[19]),
  .I1(sdpb_inst_103_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1217 (
  .O(mux_o_1217),
  .I0(sdpb_inst_104_dout[19]),
  .I1(sdpb_inst_105_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1218 (
  .O(mux_o_1218),
  .I0(sdpb_inst_106_dout[19]),
  .I1(sdpb_inst_107_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1219 (
  .O(mux_o_1219),
  .I0(sdpb_inst_108_dout[19]),
  .I1(sdpb_inst_109_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1220 (
  .O(mux_o_1220),
  .I0(sdpb_inst_110_dout[19]),
  .I1(sdpb_inst_111_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1221 (
  .O(mux_o_1221),
  .I0(sdpb_inst_112_dout[19]),
  .I1(sdpb_inst_113_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1222 (
  .O(mux_o_1222),
  .I0(sdpb_inst_114_dout[19]),
  .I1(sdpb_inst_115_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1223 (
  .O(mux_o_1223),
  .I0(sdpb_inst_116_dout[19]),
  .I1(sdpb_inst_117_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1224 (
  .O(mux_o_1224),
  .I0(sdpb_inst_118_dout[19]),
  .I1(sdpb_inst_119_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1225 (
  .O(mux_o_1225),
  .I0(sdpb_inst_120_dout[19]),
  .I1(sdpb_inst_121_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1226 (
  .O(mux_o_1226),
  .I0(sdpb_inst_122_dout[19]),
  .I1(sdpb_inst_123_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1227 (
  .O(mux_o_1227),
  .I0(sdpb_inst_124_dout[19]),
  .I1(sdpb_inst_125_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1228 (
  .O(mux_o_1228),
  .I0(sdpb_inst_126_dout[19]),
  .I1(sdpb_inst_127_dout[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1229 (
  .O(mux_o_1229),
  .I0(mux_o_1197),
  .I1(mux_o_1198),
  .S0(dff_q_4)
);
MUX2 mux_inst_1230 (
  .O(mux_o_1230),
  .I0(mux_o_1199),
  .I1(mux_o_1200),
  .S0(dff_q_4)
);
MUX2 mux_inst_1231 (
  .O(mux_o_1231),
  .I0(mux_o_1201),
  .I1(mux_o_1202),
  .S0(dff_q_4)
);
MUX2 mux_inst_1232 (
  .O(mux_o_1232),
  .I0(mux_o_1203),
  .I1(mux_o_1204),
  .S0(dff_q_4)
);
MUX2 mux_inst_1233 (
  .O(mux_o_1233),
  .I0(mux_o_1205),
  .I1(mux_o_1206),
  .S0(dff_q_4)
);
MUX2 mux_inst_1234 (
  .O(mux_o_1234),
  .I0(mux_o_1207),
  .I1(mux_o_1208),
  .S0(dff_q_4)
);
MUX2 mux_inst_1235 (
  .O(mux_o_1235),
  .I0(mux_o_1209),
  .I1(mux_o_1210),
  .S0(dff_q_4)
);
MUX2 mux_inst_1236 (
  .O(mux_o_1236),
  .I0(mux_o_1211),
  .I1(mux_o_1212),
  .S0(dff_q_4)
);
MUX2 mux_inst_1237 (
  .O(mux_o_1237),
  .I0(mux_o_1213),
  .I1(mux_o_1214),
  .S0(dff_q_4)
);
MUX2 mux_inst_1238 (
  .O(mux_o_1238),
  .I0(mux_o_1215),
  .I1(mux_o_1216),
  .S0(dff_q_4)
);
MUX2 mux_inst_1239 (
  .O(mux_o_1239),
  .I0(mux_o_1217),
  .I1(mux_o_1218),
  .S0(dff_q_4)
);
MUX2 mux_inst_1240 (
  .O(mux_o_1240),
  .I0(mux_o_1219),
  .I1(mux_o_1220),
  .S0(dff_q_4)
);
MUX2 mux_inst_1241 (
  .O(mux_o_1241),
  .I0(mux_o_1221),
  .I1(mux_o_1222),
  .S0(dff_q_4)
);
MUX2 mux_inst_1242 (
  .O(mux_o_1242),
  .I0(mux_o_1223),
  .I1(mux_o_1224),
  .S0(dff_q_4)
);
MUX2 mux_inst_1243 (
  .O(mux_o_1243),
  .I0(mux_o_1225),
  .I1(mux_o_1226),
  .S0(dff_q_4)
);
MUX2 mux_inst_1244 (
  .O(mux_o_1244),
  .I0(mux_o_1227),
  .I1(mux_o_1228),
  .S0(dff_q_4)
);
MUX2 mux_inst_1245 (
  .O(mux_o_1245),
  .I0(mux_o_1229),
  .I1(mux_o_1230),
  .S0(dff_q_3)
);
MUX2 mux_inst_1246 (
  .O(mux_o_1246),
  .I0(mux_o_1231),
  .I1(mux_o_1232),
  .S0(dff_q_3)
);
MUX2 mux_inst_1247 (
  .O(mux_o_1247),
  .I0(mux_o_1233),
  .I1(mux_o_1234),
  .S0(dff_q_3)
);
MUX2 mux_inst_1248 (
  .O(mux_o_1248),
  .I0(mux_o_1235),
  .I1(mux_o_1236),
  .S0(dff_q_3)
);
MUX2 mux_inst_1249 (
  .O(mux_o_1249),
  .I0(mux_o_1237),
  .I1(mux_o_1238),
  .S0(dff_q_3)
);
MUX2 mux_inst_1250 (
  .O(mux_o_1250),
  .I0(mux_o_1239),
  .I1(mux_o_1240),
  .S0(dff_q_3)
);
MUX2 mux_inst_1251 (
  .O(mux_o_1251),
  .I0(mux_o_1241),
  .I1(mux_o_1242),
  .S0(dff_q_3)
);
MUX2 mux_inst_1252 (
  .O(mux_o_1252),
  .I0(mux_o_1243),
  .I1(mux_o_1244),
  .S0(dff_q_3)
);
MUX2 mux_inst_1253 (
  .O(mux_o_1253),
  .I0(mux_o_1245),
  .I1(mux_o_1246),
  .S0(dff_q_2)
);
MUX2 mux_inst_1254 (
  .O(mux_o_1254),
  .I0(mux_o_1247),
  .I1(mux_o_1248),
  .S0(dff_q_2)
);
MUX2 mux_inst_1255 (
  .O(mux_o_1255),
  .I0(mux_o_1249),
  .I1(mux_o_1250),
  .S0(dff_q_2)
);
MUX2 mux_inst_1256 (
  .O(mux_o_1256),
  .I0(mux_o_1251),
  .I1(mux_o_1252),
  .S0(dff_q_2)
);
MUX2 mux_inst_1257 (
  .O(mux_o_1257),
  .I0(mux_o_1253),
  .I1(mux_o_1254),
  .S0(dff_q_1)
);
MUX2 mux_inst_1258 (
  .O(mux_o_1258),
  .I0(mux_o_1255),
  .I1(mux_o_1256),
  .S0(dff_q_1)
);
MUX2 mux_inst_1259 (
  .O(dout[19]),
  .I0(mux_o_1257),
  .I1(mux_o_1258),
  .S0(dff_q_0)
);
MUX2 mux_inst_1260 (
  .O(mux_o_1260),
  .I0(sdpb_inst_64_dout[20]),
  .I1(sdpb_inst_65_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1261 (
  .O(mux_o_1261),
  .I0(sdpb_inst_66_dout[20]),
  .I1(sdpb_inst_67_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1262 (
  .O(mux_o_1262),
  .I0(sdpb_inst_68_dout[20]),
  .I1(sdpb_inst_69_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1263 (
  .O(mux_o_1263),
  .I0(sdpb_inst_70_dout[20]),
  .I1(sdpb_inst_71_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1264 (
  .O(mux_o_1264),
  .I0(sdpb_inst_72_dout[20]),
  .I1(sdpb_inst_73_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1265 (
  .O(mux_o_1265),
  .I0(sdpb_inst_74_dout[20]),
  .I1(sdpb_inst_75_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1266 (
  .O(mux_o_1266),
  .I0(sdpb_inst_76_dout[20]),
  .I1(sdpb_inst_77_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1267 (
  .O(mux_o_1267),
  .I0(sdpb_inst_78_dout[20]),
  .I1(sdpb_inst_79_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1268 (
  .O(mux_o_1268),
  .I0(sdpb_inst_80_dout[20]),
  .I1(sdpb_inst_81_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1269 (
  .O(mux_o_1269),
  .I0(sdpb_inst_82_dout[20]),
  .I1(sdpb_inst_83_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1270 (
  .O(mux_o_1270),
  .I0(sdpb_inst_84_dout[20]),
  .I1(sdpb_inst_85_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1271 (
  .O(mux_o_1271),
  .I0(sdpb_inst_86_dout[20]),
  .I1(sdpb_inst_87_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1272 (
  .O(mux_o_1272),
  .I0(sdpb_inst_88_dout[20]),
  .I1(sdpb_inst_89_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1273 (
  .O(mux_o_1273),
  .I0(sdpb_inst_90_dout[20]),
  .I1(sdpb_inst_91_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1274 (
  .O(mux_o_1274),
  .I0(sdpb_inst_92_dout[20]),
  .I1(sdpb_inst_93_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1275 (
  .O(mux_o_1275),
  .I0(sdpb_inst_94_dout[20]),
  .I1(sdpb_inst_95_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1276 (
  .O(mux_o_1276),
  .I0(sdpb_inst_96_dout[20]),
  .I1(sdpb_inst_97_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1277 (
  .O(mux_o_1277),
  .I0(sdpb_inst_98_dout[20]),
  .I1(sdpb_inst_99_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1278 (
  .O(mux_o_1278),
  .I0(sdpb_inst_100_dout[20]),
  .I1(sdpb_inst_101_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1279 (
  .O(mux_o_1279),
  .I0(sdpb_inst_102_dout[20]),
  .I1(sdpb_inst_103_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1280 (
  .O(mux_o_1280),
  .I0(sdpb_inst_104_dout[20]),
  .I1(sdpb_inst_105_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1281 (
  .O(mux_o_1281),
  .I0(sdpb_inst_106_dout[20]),
  .I1(sdpb_inst_107_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1282 (
  .O(mux_o_1282),
  .I0(sdpb_inst_108_dout[20]),
  .I1(sdpb_inst_109_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1283 (
  .O(mux_o_1283),
  .I0(sdpb_inst_110_dout[20]),
  .I1(sdpb_inst_111_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1284 (
  .O(mux_o_1284),
  .I0(sdpb_inst_112_dout[20]),
  .I1(sdpb_inst_113_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1285 (
  .O(mux_o_1285),
  .I0(sdpb_inst_114_dout[20]),
  .I1(sdpb_inst_115_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1286 (
  .O(mux_o_1286),
  .I0(sdpb_inst_116_dout[20]),
  .I1(sdpb_inst_117_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1287 (
  .O(mux_o_1287),
  .I0(sdpb_inst_118_dout[20]),
  .I1(sdpb_inst_119_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1288 (
  .O(mux_o_1288),
  .I0(sdpb_inst_120_dout[20]),
  .I1(sdpb_inst_121_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1289 (
  .O(mux_o_1289),
  .I0(sdpb_inst_122_dout[20]),
  .I1(sdpb_inst_123_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1290 (
  .O(mux_o_1290),
  .I0(sdpb_inst_124_dout[20]),
  .I1(sdpb_inst_125_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1291 (
  .O(mux_o_1291),
  .I0(sdpb_inst_126_dout[20]),
  .I1(sdpb_inst_127_dout[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1292 (
  .O(mux_o_1292),
  .I0(mux_o_1260),
  .I1(mux_o_1261),
  .S0(dff_q_4)
);
MUX2 mux_inst_1293 (
  .O(mux_o_1293),
  .I0(mux_o_1262),
  .I1(mux_o_1263),
  .S0(dff_q_4)
);
MUX2 mux_inst_1294 (
  .O(mux_o_1294),
  .I0(mux_o_1264),
  .I1(mux_o_1265),
  .S0(dff_q_4)
);
MUX2 mux_inst_1295 (
  .O(mux_o_1295),
  .I0(mux_o_1266),
  .I1(mux_o_1267),
  .S0(dff_q_4)
);
MUX2 mux_inst_1296 (
  .O(mux_o_1296),
  .I0(mux_o_1268),
  .I1(mux_o_1269),
  .S0(dff_q_4)
);
MUX2 mux_inst_1297 (
  .O(mux_o_1297),
  .I0(mux_o_1270),
  .I1(mux_o_1271),
  .S0(dff_q_4)
);
MUX2 mux_inst_1298 (
  .O(mux_o_1298),
  .I0(mux_o_1272),
  .I1(mux_o_1273),
  .S0(dff_q_4)
);
MUX2 mux_inst_1299 (
  .O(mux_o_1299),
  .I0(mux_o_1274),
  .I1(mux_o_1275),
  .S0(dff_q_4)
);
MUX2 mux_inst_1300 (
  .O(mux_o_1300),
  .I0(mux_o_1276),
  .I1(mux_o_1277),
  .S0(dff_q_4)
);
MUX2 mux_inst_1301 (
  .O(mux_o_1301),
  .I0(mux_o_1278),
  .I1(mux_o_1279),
  .S0(dff_q_4)
);
MUX2 mux_inst_1302 (
  .O(mux_o_1302),
  .I0(mux_o_1280),
  .I1(mux_o_1281),
  .S0(dff_q_4)
);
MUX2 mux_inst_1303 (
  .O(mux_o_1303),
  .I0(mux_o_1282),
  .I1(mux_o_1283),
  .S0(dff_q_4)
);
MUX2 mux_inst_1304 (
  .O(mux_o_1304),
  .I0(mux_o_1284),
  .I1(mux_o_1285),
  .S0(dff_q_4)
);
MUX2 mux_inst_1305 (
  .O(mux_o_1305),
  .I0(mux_o_1286),
  .I1(mux_o_1287),
  .S0(dff_q_4)
);
MUX2 mux_inst_1306 (
  .O(mux_o_1306),
  .I0(mux_o_1288),
  .I1(mux_o_1289),
  .S0(dff_q_4)
);
MUX2 mux_inst_1307 (
  .O(mux_o_1307),
  .I0(mux_o_1290),
  .I1(mux_o_1291),
  .S0(dff_q_4)
);
MUX2 mux_inst_1308 (
  .O(mux_o_1308),
  .I0(mux_o_1292),
  .I1(mux_o_1293),
  .S0(dff_q_3)
);
MUX2 mux_inst_1309 (
  .O(mux_o_1309),
  .I0(mux_o_1294),
  .I1(mux_o_1295),
  .S0(dff_q_3)
);
MUX2 mux_inst_1310 (
  .O(mux_o_1310),
  .I0(mux_o_1296),
  .I1(mux_o_1297),
  .S0(dff_q_3)
);
MUX2 mux_inst_1311 (
  .O(mux_o_1311),
  .I0(mux_o_1298),
  .I1(mux_o_1299),
  .S0(dff_q_3)
);
MUX2 mux_inst_1312 (
  .O(mux_o_1312),
  .I0(mux_o_1300),
  .I1(mux_o_1301),
  .S0(dff_q_3)
);
MUX2 mux_inst_1313 (
  .O(mux_o_1313),
  .I0(mux_o_1302),
  .I1(mux_o_1303),
  .S0(dff_q_3)
);
MUX2 mux_inst_1314 (
  .O(mux_o_1314),
  .I0(mux_o_1304),
  .I1(mux_o_1305),
  .S0(dff_q_3)
);
MUX2 mux_inst_1315 (
  .O(mux_o_1315),
  .I0(mux_o_1306),
  .I1(mux_o_1307),
  .S0(dff_q_3)
);
MUX2 mux_inst_1316 (
  .O(mux_o_1316),
  .I0(mux_o_1308),
  .I1(mux_o_1309),
  .S0(dff_q_2)
);
MUX2 mux_inst_1317 (
  .O(mux_o_1317),
  .I0(mux_o_1310),
  .I1(mux_o_1311),
  .S0(dff_q_2)
);
MUX2 mux_inst_1318 (
  .O(mux_o_1318),
  .I0(mux_o_1312),
  .I1(mux_o_1313),
  .S0(dff_q_2)
);
MUX2 mux_inst_1319 (
  .O(mux_o_1319),
  .I0(mux_o_1314),
  .I1(mux_o_1315),
  .S0(dff_q_2)
);
MUX2 mux_inst_1320 (
  .O(mux_o_1320),
  .I0(mux_o_1316),
  .I1(mux_o_1317),
  .S0(dff_q_1)
);
MUX2 mux_inst_1321 (
  .O(mux_o_1321),
  .I0(mux_o_1318),
  .I1(mux_o_1319),
  .S0(dff_q_1)
);
MUX2 mux_inst_1322 (
  .O(dout[20]),
  .I0(mux_o_1320),
  .I1(mux_o_1321),
  .S0(dff_q_0)
);
MUX2 mux_inst_1323 (
  .O(mux_o_1323),
  .I0(sdpb_inst_64_dout[21]),
  .I1(sdpb_inst_65_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1324 (
  .O(mux_o_1324),
  .I0(sdpb_inst_66_dout[21]),
  .I1(sdpb_inst_67_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1325 (
  .O(mux_o_1325),
  .I0(sdpb_inst_68_dout[21]),
  .I1(sdpb_inst_69_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1326 (
  .O(mux_o_1326),
  .I0(sdpb_inst_70_dout[21]),
  .I1(sdpb_inst_71_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1327 (
  .O(mux_o_1327),
  .I0(sdpb_inst_72_dout[21]),
  .I1(sdpb_inst_73_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1328 (
  .O(mux_o_1328),
  .I0(sdpb_inst_74_dout[21]),
  .I1(sdpb_inst_75_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1329 (
  .O(mux_o_1329),
  .I0(sdpb_inst_76_dout[21]),
  .I1(sdpb_inst_77_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1330 (
  .O(mux_o_1330),
  .I0(sdpb_inst_78_dout[21]),
  .I1(sdpb_inst_79_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1331 (
  .O(mux_o_1331),
  .I0(sdpb_inst_80_dout[21]),
  .I1(sdpb_inst_81_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1332 (
  .O(mux_o_1332),
  .I0(sdpb_inst_82_dout[21]),
  .I1(sdpb_inst_83_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1333 (
  .O(mux_o_1333),
  .I0(sdpb_inst_84_dout[21]),
  .I1(sdpb_inst_85_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1334 (
  .O(mux_o_1334),
  .I0(sdpb_inst_86_dout[21]),
  .I1(sdpb_inst_87_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1335 (
  .O(mux_o_1335),
  .I0(sdpb_inst_88_dout[21]),
  .I1(sdpb_inst_89_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1336 (
  .O(mux_o_1336),
  .I0(sdpb_inst_90_dout[21]),
  .I1(sdpb_inst_91_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1337 (
  .O(mux_o_1337),
  .I0(sdpb_inst_92_dout[21]),
  .I1(sdpb_inst_93_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1338 (
  .O(mux_o_1338),
  .I0(sdpb_inst_94_dout[21]),
  .I1(sdpb_inst_95_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1339 (
  .O(mux_o_1339),
  .I0(sdpb_inst_96_dout[21]),
  .I1(sdpb_inst_97_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1340 (
  .O(mux_o_1340),
  .I0(sdpb_inst_98_dout[21]),
  .I1(sdpb_inst_99_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1341 (
  .O(mux_o_1341),
  .I0(sdpb_inst_100_dout[21]),
  .I1(sdpb_inst_101_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1342 (
  .O(mux_o_1342),
  .I0(sdpb_inst_102_dout[21]),
  .I1(sdpb_inst_103_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1343 (
  .O(mux_o_1343),
  .I0(sdpb_inst_104_dout[21]),
  .I1(sdpb_inst_105_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1344 (
  .O(mux_o_1344),
  .I0(sdpb_inst_106_dout[21]),
  .I1(sdpb_inst_107_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1345 (
  .O(mux_o_1345),
  .I0(sdpb_inst_108_dout[21]),
  .I1(sdpb_inst_109_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1346 (
  .O(mux_o_1346),
  .I0(sdpb_inst_110_dout[21]),
  .I1(sdpb_inst_111_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1347 (
  .O(mux_o_1347),
  .I0(sdpb_inst_112_dout[21]),
  .I1(sdpb_inst_113_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1348 (
  .O(mux_o_1348),
  .I0(sdpb_inst_114_dout[21]),
  .I1(sdpb_inst_115_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1349 (
  .O(mux_o_1349),
  .I0(sdpb_inst_116_dout[21]),
  .I1(sdpb_inst_117_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1350 (
  .O(mux_o_1350),
  .I0(sdpb_inst_118_dout[21]),
  .I1(sdpb_inst_119_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1351 (
  .O(mux_o_1351),
  .I0(sdpb_inst_120_dout[21]),
  .I1(sdpb_inst_121_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1352 (
  .O(mux_o_1352),
  .I0(sdpb_inst_122_dout[21]),
  .I1(sdpb_inst_123_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1353 (
  .O(mux_o_1353),
  .I0(sdpb_inst_124_dout[21]),
  .I1(sdpb_inst_125_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1354 (
  .O(mux_o_1354),
  .I0(sdpb_inst_126_dout[21]),
  .I1(sdpb_inst_127_dout[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1355 (
  .O(mux_o_1355),
  .I0(mux_o_1323),
  .I1(mux_o_1324),
  .S0(dff_q_4)
);
MUX2 mux_inst_1356 (
  .O(mux_o_1356),
  .I0(mux_o_1325),
  .I1(mux_o_1326),
  .S0(dff_q_4)
);
MUX2 mux_inst_1357 (
  .O(mux_o_1357),
  .I0(mux_o_1327),
  .I1(mux_o_1328),
  .S0(dff_q_4)
);
MUX2 mux_inst_1358 (
  .O(mux_o_1358),
  .I0(mux_o_1329),
  .I1(mux_o_1330),
  .S0(dff_q_4)
);
MUX2 mux_inst_1359 (
  .O(mux_o_1359),
  .I0(mux_o_1331),
  .I1(mux_o_1332),
  .S0(dff_q_4)
);
MUX2 mux_inst_1360 (
  .O(mux_o_1360),
  .I0(mux_o_1333),
  .I1(mux_o_1334),
  .S0(dff_q_4)
);
MUX2 mux_inst_1361 (
  .O(mux_o_1361),
  .I0(mux_o_1335),
  .I1(mux_o_1336),
  .S0(dff_q_4)
);
MUX2 mux_inst_1362 (
  .O(mux_o_1362),
  .I0(mux_o_1337),
  .I1(mux_o_1338),
  .S0(dff_q_4)
);
MUX2 mux_inst_1363 (
  .O(mux_o_1363),
  .I0(mux_o_1339),
  .I1(mux_o_1340),
  .S0(dff_q_4)
);
MUX2 mux_inst_1364 (
  .O(mux_o_1364),
  .I0(mux_o_1341),
  .I1(mux_o_1342),
  .S0(dff_q_4)
);
MUX2 mux_inst_1365 (
  .O(mux_o_1365),
  .I0(mux_o_1343),
  .I1(mux_o_1344),
  .S0(dff_q_4)
);
MUX2 mux_inst_1366 (
  .O(mux_o_1366),
  .I0(mux_o_1345),
  .I1(mux_o_1346),
  .S0(dff_q_4)
);
MUX2 mux_inst_1367 (
  .O(mux_o_1367),
  .I0(mux_o_1347),
  .I1(mux_o_1348),
  .S0(dff_q_4)
);
MUX2 mux_inst_1368 (
  .O(mux_o_1368),
  .I0(mux_o_1349),
  .I1(mux_o_1350),
  .S0(dff_q_4)
);
MUX2 mux_inst_1369 (
  .O(mux_o_1369),
  .I0(mux_o_1351),
  .I1(mux_o_1352),
  .S0(dff_q_4)
);
MUX2 mux_inst_1370 (
  .O(mux_o_1370),
  .I0(mux_o_1353),
  .I1(mux_o_1354),
  .S0(dff_q_4)
);
MUX2 mux_inst_1371 (
  .O(mux_o_1371),
  .I0(mux_o_1355),
  .I1(mux_o_1356),
  .S0(dff_q_3)
);
MUX2 mux_inst_1372 (
  .O(mux_o_1372),
  .I0(mux_o_1357),
  .I1(mux_o_1358),
  .S0(dff_q_3)
);
MUX2 mux_inst_1373 (
  .O(mux_o_1373),
  .I0(mux_o_1359),
  .I1(mux_o_1360),
  .S0(dff_q_3)
);
MUX2 mux_inst_1374 (
  .O(mux_o_1374),
  .I0(mux_o_1361),
  .I1(mux_o_1362),
  .S0(dff_q_3)
);
MUX2 mux_inst_1375 (
  .O(mux_o_1375),
  .I0(mux_o_1363),
  .I1(mux_o_1364),
  .S0(dff_q_3)
);
MUX2 mux_inst_1376 (
  .O(mux_o_1376),
  .I0(mux_o_1365),
  .I1(mux_o_1366),
  .S0(dff_q_3)
);
MUX2 mux_inst_1377 (
  .O(mux_o_1377),
  .I0(mux_o_1367),
  .I1(mux_o_1368),
  .S0(dff_q_3)
);
MUX2 mux_inst_1378 (
  .O(mux_o_1378),
  .I0(mux_o_1369),
  .I1(mux_o_1370),
  .S0(dff_q_3)
);
MUX2 mux_inst_1379 (
  .O(mux_o_1379),
  .I0(mux_o_1371),
  .I1(mux_o_1372),
  .S0(dff_q_2)
);
MUX2 mux_inst_1380 (
  .O(mux_o_1380),
  .I0(mux_o_1373),
  .I1(mux_o_1374),
  .S0(dff_q_2)
);
MUX2 mux_inst_1381 (
  .O(mux_o_1381),
  .I0(mux_o_1375),
  .I1(mux_o_1376),
  .S0(dff_q_2)
);
MUX2 mux_inst_1382 (
  .O(mux_o_1382),
  .I0(mux_o_1377),
  .I1(mux_o_1378),
  .S0(dff_q_2)
);
MUX2 mux_inst_1383 (
  .O(mux_o_1383),
  .I0(mux_o_1379),
  .I1(mux_o_1380),
  .S0(dff_q_1)
);
MUX2 mux_inst_1384 (
  .O(mux_o_1384),
  .I0(mux_o_1381),
  .I1(mux_o_1382),
  .S0(dff_q_1)
);
MUX2 mux_inst_1385 (
  .O(dout[21]),
  .I0(mux_o_1383),
  .I1(mux_o_1384),
  .S0(dff_q_0)
);
MUX2 mux_inst_1386 (
  .O(mux_o_1386),
  .I0(sdpb_inst_64_dout[22]),
  .I1(sdpb_inst_65_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1387 (
  .O(mux_o_1387),
  .I0(sdpb_inst_66_dout[22]),
  .I1(sdpb_inst_67_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1388 (
  .O(mux_o_1388),
  .I0(sdpb_inst_68_dout[22]),
  .I1(sdpb_inst_69_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1389 (
  .O(mux_o_1389),
  .I0(sdpb_inst_70_dout[22]),
  .I1(sdpb_inst_71_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1390 (
  .O(mux_o_1390),
  .I0(sdpb_inst_72_dout[22]),
  .I1(sdpb_inst_73_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1391 (
  .O(mux_o_1391),
  .I0(sdpb_inst_74_dout[22]),
  .I1(sdpb_inst_75_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1392 (
  .O(mux_o_1392),
  .I0(sdpb_inst_76_dout[22]),
  .I1(sdpb_inst_77_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1393 (
  .O(mux_o_1393),
  .I0(sdpb_inst_78_dout[22]),
  .I1(sdpb_inst_79_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1394 (
  .O(mux_o_1394),
  .I0(sdpb_inst_80_dout[22]),
  .I1(sdpb_inst_81_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1395 (
  .O(mux_o_1395),
  .I0(sdpb_inst_82_dout[22]),
  .I1(sdpb_inst_83_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1396 (
  .O(mux_o_1396),
  .I0(sdpb_inst_84_dout[22]),
  .I1(sdpb_inst_85_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1397 (
  .O(mux_o_1397),
  .I0(sdpb_inst_86_dout[22]),
  .I1(sdpb_inst_87_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1398 (
  .O(mux_o_1398),
  .I0(sdpb_inst_88_dout[22]),
  .I1(sdpb_inst_89_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1399 (
  .O(mux_o_1399),
  .I0(sdpb_inst_90_dout[22]),
  .I1(sdpb_inst_91_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1400 (
  .O(mux_o_1400),
  .I0(sdpb_inst_92_dout[22]),
  .I1(sdpb_inst_93_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1401 (
  .O(mux_o_1401),
  .I0(sdpb_inst_94_dout[22]),
  .I1(sdpb_inst_95_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1402 (
  .O(mux_o_1402),
  .I0(sdpb_inst_96_dout[22]),
  .I1(sdpb_inst_97_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1403 (
  .O(mux_o_1403),
  .I0(sdpb_inst_98_dout[22]),
  .I1(sdpb_inst_99_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1404 (
  .O(mux_o_1404),
  .I0(sdpb_inst_100_dout[22]),
  .I1(sdpb_inst_101_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1405 (
  .O(mux_o_1405),
  .I0(sdpb_inst_102_dout[22]),
  .I1(sdpb_inst_103_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1406 (
  .O(mux_o_1406),
  .I0(sdpb_inst_104_dout[22]),
  .I1(sdpb_inst_105_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1407 (
  .O(mux_o_1407),
  .I0(sdpb_inst_106_dout[22]),
  .I1(sdpb_inst_107_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1408 (
  .O(mux_o_1408),
  .I0(sdpb_inst_108_dout[22]),
  .I1(sdpb_inst_109_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1409 (
  .O(mux_o_1409),
  .I0(sdpb_inst_110_dout[22]),
  .I1(sdpb_inst_111_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1410 (
  .O(mux_o_1410),
  .I0(sdpb_inst_112_dout[22]),
  .I1(sdpb_inst_113_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1411 (
  .O(mux_o_1411),
  .I0(sdpb_inst_114_dout[22]),
  .I1(sdpb_inst_115_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1412 (
  .O(mux_o_1412),
  .I0(sdpb_inst_116_dout[22]),
  .I1(sdpb_inst_117_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1413 (
  .O(mux_o_1413),
  .I0(sdpb_inst_118_dout[22]),
  .I1(sdpb_inst_119_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1414 (
  .O(mux_o_1414),
  .I0(sdpb_inst_120_dout[22]),
  .I1(sdpb_inst_121_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1415 (
  .O(mux_o_1415),
  .I0(sdpb_inst_122_dout[22]),
  .I1(sdpb_inst_123_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1416 (
  .O(mux_o_1416),
  .I0(sdpb_inst_124_dout[22]),
  .I1(sdpb_inst_125_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1417 (
  .O(mux_o_1417),
  .I0(sdpb_inst_126_dout[22]),
  .I1(sdpb_inst_127_dout[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1418 (
  .O(mux_o_1418),
  .I0(mux_o_1386),
  .I1(mux_o_1387),
  .S0(dff_q_4)
);
MUX2 mux_inst_1419 (
  .O(mux_o_1419),
  .I0(mux_o_1388),
  .I1(mux_o_1389),
  .S0(dff_q_4)
);
MUX2 mux_inst_1420 (
  .O(mux_o_1420),
  .I0(mux_o_1390),
  .I1(mux_o_1391),
  .S0(dff_q_4)
);
MUX2 mux_inst_1421 (
  .O(mux_o_1421),
  .I0(mux_o_1392),
  .I1(mux_o_1393),
  .S0(dff_q_4)
);
MUX2 mux_inst_1422 (
  .O(mux_o_1422),
  .I0(mux_o_1394),
  .I1(mux_o_1395),
  .S0(dff_q_4)
);
MUX2 mux_inst_1423 (
  .O(mux_o_1423),
  .I0(mux_o_1396),
  .I1(mux_o_1397),
  .S0(dff_q_4)
);
MUX2 mux_inst_1424 (
  .O(mux_o_1424),
  .I0(mux_o_1398),
  .I1(mux_o_1399),
  .S0(dff_q_4)
);
MUX2 mux_inst_1425 (
  .O(mux_o_1425),
  .I0(mux_o_1400),
  .I1(mux_o_1401),
  .S0(dff_q_4)
);
MUX2 mux_inst_1426 (
  .O(mux_o_1426),
  .I0(mux_o_1402),
  .I1(mux_o_1403),
  .S0(dff_q_4)
);
MUX2 mux_inst_1427 (
  .O(mux_o_1427),
  .I0(mux_o_1404),
  .I1(mux_o_1405),
  .S0(dff_q_4)
);
MUX2 mux_inst_1428 (
  .O(mux_o_1428),
  .I0(mux_o_1406),
  .I1(mux_o_1407),
  .S0(dff_q_4)
);
MUX2 mux_inst_1429 (
  .O(mux_o_1429),
  .I0(mux_o_1408),
  .I1(mux_o_1409),
  .S0(dff_q_4)
);
MUX2 mux_inst_1430 (
  .O(mux_o_1430),
  .I0(mux_o_1410),
  .I1(mux_o_1411),
  .S0(dff_q_4)
);
MUX2 mux_inst_1431 (
  .O(mux_o_1431),
  .I0(mux_o_1412),
  .I1(mux_o_1413),
  .S0(dff_q_4)
);
MUX2 mux_inst_1432 (
  .O(mux_o_1432),
  .I0(mux_o_1414),
  .I1(mux_o_1415),
  .S0(dff_q_4)
);
MUX2 mux_inst_1433 (
  .O(mux_o_1433),
  .I0(mux_o_1416),
  .I1(mux_o_1417),
  .S0(dff_q_4)
);
MUX2 mux_inst_1434 (
  .O(mux_o_1434),
  .I0(mux_o_1418),
  .I1(mux_o_1419),
  .S0(dff_q_3)
);
MUX2 mux_inst_1435 (
  .O(mux_o_1435),
  .I0(mux_o_1420),
  .I1(mux_o_1421),
  .S0(dff_q_3)
);
MUX2 mux_inst_1436 (
  .O(mux_o_1436),
  .I0(mux_o_1422),
  .I1(mux_o_1423),
  .S0(dff_q_3)
);
MUX2 mux_inst_1437 (
  .O(mux_o_1437),
  .I0(mux_o_1424),
  .I1(mux_o_1425),
  .S0(dff_q_3)
);
MUX2 mux_inst_1438 (
  .O(mux_o_1438),
  .I0(mux_o_1426),
  .I1(mux_o_1427),
  .S0(dff_q_3)
);
MUX2 mux_inst_1439 (
  .O(mux_o_1439),
  .I0(mux_o_1428),
  .I1(mux_o_1429),
  .S0(dff_q_3)
);
MUX2 mux_inst_1440 (
  .O(mux_o_1440),
  .I0(mux_o_1430),
  .I1(mux_o_1431),
  .S0(dff_q_3)
);
MUX2 mux_inst_1441 (
  .O(mux_o_1441),
  .I0(mux_o_1432),
  .I1(mux_o_1433),
  .S0(dff_q_3)
);
MUX2 mux_inst_1442 (
  .O(mux_o_1442),
  .I0(mux_o_1434),
  .I1(mux_o_1435),
  .S0(dff_q_2)
);
MUX2 mux_inst_1443 (
  .O(mux_o_1443),
  .I0(mux_o_1436),
  .I1(mux_o_1437),
  .S0(dff_q_2)
);
MUX2 mux_inst_1444 (
  .O(mux_o_1444),
  .I0(mux_o_1438),
  .I1(mux_o_1439),
  .S0(dff_q_2)
);
MUX2 mux_inst_1445 (
  .O(mux_o_1445),
  .I0(mux_o_1440),
  .I1(mux_o_1441),
  .S0(dff_q_2)
);
MUX2 mux_inst_1446 (
  .O(mux_o_1446),
  .I0(mux_o_1442),
  .I1(mux_o_1443),
  .S0(dff_q_1)
);
MUX2 mux_inst_1447 (
  .O(mux_o_1447),
  .I0(mux_o_1444),
  .I1(mux_o_1445),
  .S0(dff_q_1)
);
MUX2 mux_inst_1448 (
  .O(dout[22]),
  .I0(mux_o_1446),
  .I1(mux_o_1447),
  .S0(dff_q_0)
);
MUX2 mux_inst_1449 (
  .O(mux_o_1449),
  .I0(sdpb_inst_64_dout[23]),
  .I1(sdpb_inst_65_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1450 (
  .O(mux_o_1450),
  .I0(sdpb_inst_66_dout[23]),
  .I1(sdpb_inst_67_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1451 (
  .O(mux_o_1451),
  .I0(sdpb_inst_68_dout[23]),
  .I1(sdpb_inst_69_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1452 (
  .O(mux_o_1452),
  .I0(sdpb_inst_70_dout[23]),
  .I1(sdpb_inst_71_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1453 (
  .O(mux_o_1453),
  .I0(sdpb_inst_72_dout[23]),
  .I1(sdpb_inst_73_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1454 (
  .O(mux_o_1454),
  .I0(sdpb_inst_74_dout[23]),
  .I1(sdpb_inst_75_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1455 (
  .O(mux_o_1455),
  .I0(sdpb_inst_76_dout[23]),
  .I1(sdpb_inst_77_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1456 (
  .O(mux_o_1456),
  .I0(sdpb_inst_78_dout[23]),
  .I1(sdpb_inst_79_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1457 (
  .O(mux_o_1457),
  .I0(sdpb_inst_80_dout[23]),
  .I1(sdpb_inst_81_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1458 (
  .O(mux_o_1458),
  .I0(sdpb_inst_82_dout[23]),
  .I1(sdpb_inst_83_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1459 (
  .O(mux_o_1459),
  .I0(sdpb_inst_84_dout[23]),
  .I1(sdpb_inst_85_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1460 (
  .O(mux_o_1460),
  .I0(sdpb_inst_86_dout[23]),
  .I1(sdpb_inst_87_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1461 (
  .O(mux_o_1461),
  .I0(sdpb_inst_88_dout[23]),
  .I1(sdpb_inst_89_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1462 (
  .O(mux_o_1462),
  .I0(sdpb_inst_90_dout[23]),
  .I1(sdpb_inst_91_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1463 (
  .O(mux_o_1463),
  .I0(sdpb_inst_92_dout[23]),
  .I1(sdpb_inst_93_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1464 (
  .O(mux_o_1464),
  .I0(sdpb_inst_94_dout[23]),
  .I1(sdpb_inst_95_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1465 (
  .O(mux_o_1465),
  .I0(sdpb_inst_96_dout[23]),
  .I1(sdpb_inst_97_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1466 (
  .O(mux_o_1466),
  .I0(sdpb_inst_98_dout[23]),
  .I1(sdpb_inst_99_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1467 (
  .O(mux_o_1467),
  .I0(sdpb_inst_100_dout[23]),
  .I1(sdpb_inst_101_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1468 (
  .O(mux_o_1468),
  .I0(sdpb_inst_102_dout[23]),
  .I1(sdpb_inst_103_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1469 (
  .O(mux_o_1469),
  .I0(sdpb_inst_104_dout[23]),
  .I1(sdpb_inst_105_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1470 (
  .O(mux_o_1470),
  .I0(sdpb_inst_106_dout[23]),
  .I1(sdpb_inst_107_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1471 (
  .O(mux_o_1471),
  .I0(sdpb_inst_108_dout[23]),
  .I1(sdpb_inst_109_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1472 (
  .O(mux_o_1472),
  .I0(sdpb_inst_110_dout[23]),
  .I1(sdpb_inst_111_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1473 (
  .O(mux_o_1473),
  .I0(sdpb_inst_112_dout[23]),
  .I1(sdpb_inst_113_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1474 (
  .O(mux_o_1474),
  .I0(sdpb_inst_114_dout[23]),
  .I1(sdpb_inst_115_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1475 (
  .O(mux_o_1475),
  .I0(sdpb_inst_116_dout[23]),
  .I1(sdpb_inst_117_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1476 (
  .O(mux_o_1476),
  .I0(sdpb_inst_118_dout[23]),
  .I1(sdpb_inst_119_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1477 (
  .O(mux_o_1477),
  .I0(sdpb_inst_120_dout[23]),
  .I1(sdpb_inst_121_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1478 (
  .O(mux_o_1478),
  .I0(sdpb_inst_122_dout[23]),
  .I1(sdpb_inst_123_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1479 (
  .O(mux_o_1479),
  .I0(sdpb_inst_124_dout[23]),
  .I1(sdpb_inst_125_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1480 (
  .O(mux_o_1480),
  .I0(sdpb_inst_126_dout[23]),
  .I1(sdpb_inst_127_dout[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1481 (
  .O(mux_o_1481),
  .I0(mux_o_1449),
  .I1(mux_o_1450),
  .S0(dff_q_4)
);
MUX2 mux_inst_1482 (
  .O(mux_o_1482),
  .I0(mux_o_1451),
  .I1(mux_o_1452),
  .S0(dff_q_4)
);
MUX2 mux_inst_1483 (
  .O(mux_o_1483),
  .I0(mux_o_1453),
  .I1(mux_o_1454),
  .S0(dff_q_4)
);
MUX2 mux_inst_1484 (
  .O(mux_o_1484),
  .I0(mux_o_1455),
  .I1(mux_o_1456),
  .S0(dff_q_4)
);
MUX2 mux_inst_1485 (
  .O(mux_o_1485),
  .I0(mux_o_1457),
  .I1(mux_o_1458),
  .S0(dff_q_4)
);
MUX2 mux_inst_1486 (
  .O(mux_o_1486),
  .I0(mux_o_1459),
  .I1(mux_o_1460),
  .S0(dff_q_4)
);
MUX2 mux_inst_1487 (
  .O(mux_o_1487),
  .I0(mux_o_1461),
  .I1(mux_o_1462),
  .S0(dff_q_4)
);
MUX2 mux_inst_1488 (
  .O(mux_o_1488),
  .I0(mux_o_1463),
  .I1(mux_o_1464),
  .S0(dff_q_4)
);
MUX2 mux_inst_1489 (
  .O(mux_o_1489),
  .I0(mux_o_1465),
  .I1(mux_o_1466),
  .S0(dff_q_4)
);
MUX2 mux_inst_1490 (
  .O(mux_o_1490),
  .I0(mux_o_1467),
  .I1(mux_o_1468),
  .S0(dff_q_4)
);
MUX2 mux_inst_1491 (
  .O(mux_o_1491),
  .I0(mux_o_1469),
  .I1(mux_o_1470),
  .S0(dff_q_4)
);
MUX2 mux_inst_1492 (
  .O(mux_o_1492),
  .I0(mux_o_1471),
  .I1(mux_o_1472),
  .S0(dff_q_4)
);
MUX2 mux_inst_1493 (
  .O(mux_o_1493),
  .I0(mux_o_1473),
  .I1(mux_o_1474),
  .S0(dff_q_4)
);
MUX2 mux_inst_1494 (
  .O(mux_o_1494),
  .I0(mux_o_1475),
  .I1(mux_o_1476),
  .S0(dff_q_4)
);
MUX2 mux_inst_1495 (
  .O(mux_o_1495),
  .I0(mux_o_1477),
  .I1(mux_o_1478),
  .S0(dff_q_4)
);
MUX2 mux_inst_1496 (
  .O(mux_o_1496),
  .I0(mux_o_1479),
  .I1(mux_o_1480),
  .S0(dff_q_4)
);
MUX2 mux_inst_1497 (
  .O(mux_o_1497),
  .I0(mux_o_1481),
  .I1(mux_o_1482),
  .S0(dff_q_3)
);
MUX2 mux_inst_1498 (
  .O(mux_o_1498),
  .I0(mux_o_1483),
  .I1(mux_o_1484),
  .S0(dff_q_3)
);
MUX2 mux_inst_1499 (
  .O(mux_o_1499),
  .I0(mux_o_1485),
  .I1(mux_o_1486),
  .S0(dff_q_3)
);
MUX2 mux_inst_1500 (
  .O(mux_o_1500),
  .I0(mux_o_1487),
  .I1(mux_o_1488),
  .S0(dff_q_3)
);
MUX2 mux_inst_1501 (
  .O(mux_o_1501),
  .I0(mux_o_1489),
  .I1(mux_o_1490),
  .S0(dff_q_3)
);
MUX2 mux_inst_1502 (
  .O(mux_o_1502),
  .I0(mux_o_1491),
  .I1(mux_o_1492),
  .S0(dff_q_3)
);
MUX2 mux_inst_1503 (
  .O(mux_o_1503),
  .I0(mux_o_1493),
  .I1(mux_o_1494),
  .S0(dff_q_3)
);
MUX2 mux_inst_1504 (
  .O(mux_o_1504),
  .I0(mux_o_1495),
  .I1(mux_o_1496),
  .S0(dff_q_3)
);
MUX2 mux_inst_1505 (
  .O(mux_o_1505),
  .I0(mux_o_1497),
  .I1(mux_o_1498),
  .S0(dff_q_2)
);
MUX2 mux_inst_1506 (
  .O(mux_o_1506),
  .I0(mux_o_1499),
  .I1(mux_o_1500),
  .S0(dff_q_2)
);
MUX2 mux_inst_1507 (
  .O(mux_o_1507),
  .I0(mux_o_1501),
  .I1(mux_o_1502),
  .S0(dff_q_2)
);
MUX2 mux_inst_1508 (
  .O(mux_o_1508),
  .I0(mux_o_1503),
  .I1(mux_o_1504),
  .S0(dff_q_2)
);
MUX2 mux_inst_1509 (
  .O(mux_o_1509),
  .I0(mux_o_1505),
  .I1(mux_o_1506),
  .S0(dff_q_1)
);
MUX2 mux_inst_1510 (
  .O(mux_o_1510),
  .I0(mux_o_1507),
  .I1(mux_o_1508),
  .S0(dff_q_1)
);
MUX2 mux_inst_1511 (
  .O(dout[23]),
  .I0(mux_o_1509),
  .I1(mux_o_1510),
  .S0(dff_q_0)
);
MUX2 mux_inst_1512 (
  .O(mux_o_1512),
  .I0(sdpb_inst_64_dout[24]),
  .I1(sdpb_inst_65_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1513 (
  .O(mux_o_1513),
  .I0(sdpb_inst_66_dout[24]),
  .I1(sdpb_inst_67_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1514 (
  .O(mux_o_1514),
  .I0(sdpb_inst_68_dout[24]),
  .I1(sdpb_inst_69_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1515 (
  .O(mux_o_1515),
  .I0(sdpb_inst_70_dout[24]),
  .I1(sdpb_inst_71_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1516 (
  .O(mux_o_1516),
  .I0(sdpb_inst_72_dout[24]),
  .I1(sdpb_inst_73_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1517 (
  .O(mux_o_1517),
  .I0(sdpb_inst_74_dout[24]),
  .I1(sdpb_inst_75_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1518 (
  .O(mux_o_1518),
  .I0(sdpb_inst_76_dout[24]),
  .I1(sdpb_inst_77_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1519 (
  .O(mux_o_1519),
  .I0(sdpb_inst_78_dout[24]),
  .I1(sdpb_inst_79_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1520 (
  .O(mux_o_1520),
  .I0(sdpb_inst_80_dout[24]),
  .I1(sdpb_inst_81_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1521 (
  .O(mux_o_1521),
  .I0(sdpb_inst_82_dout[24]),
  .I1(sdpb_inst_83_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1522 (
  .O(mux_o_1522),
  .I0(sdpb_inst_84_dout[24]),
  .I1(sdpb_inst_85_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1523 (
  .O(mux_o_1523),
  .I0(sdpb_inst_86_dout[24]),
  .I1(sdpb_inst_87_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1524 (
  .O(mux_o_1524),
  .I0(sdpb_inst_88_dout[24]),
  .I1(sdpb_inst_89_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1525 (
  .O(mux_o_1525),
  .I0(sdpb_inst_90_dout[24]),
  .I1(sdpb_inst_91_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1526 (
  .O(mux_o_1526),
  .I0(sdpb_inst_92_dout[24]),
  .I1(sdpb_inst_93_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1527 (
  .O(mux_o_1527),
  .I0(sdpb_inst_94_dout[24]),
  .I1(sdpb_inst_95_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1528 (
  .O(mux_o_1528),
  .I0(sdpb_inst_96_dout[24]),
  .I1(sdpb_inst_97_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1529 (
  .O(mux_o_1529),
  .I0(sdpb_inst_98_dout[24]),
  .I1(sdpb_inst_99_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1530 (
  .O(mux_o_1530),
  .I0(sdpb_inst_100_dout[24]),
  .I1(sdpb_inst_101_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1531 (
  .O(mux_o_1531),
  .I0(sdpb_inst_102_dout[24]),
  .I1(sdpb_inst_103_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1532 (
  .O(mux_o_1532),
  .I0(sdpb_inst_104_dout[24]),
  .I1(sdpb_inst_105_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1533 (
  .O(mux_o_1533),
  .I0(sdpb_inst_106_dout[24]),
  .I1(sdpb_inst_107_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1534 (
  .O(mux_o_1534),
  .I0(sdpb_inst_108_dout[24]),
  .I1(sdpb_inst_109_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1535 (
  .O(mux_o_1535),
  .I0(sdpb_inst_110_dout[24]),
  .I1(sdpb_inst_111_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1536 (
  .O(mux_o_1536),
  .I0(sdpb_inst_112_dout[24]),
  .I1(sdpb_inst_113_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1537 (
  .O(mux_o_1537),
  .I0(sdpb_inst_114_dout[24]),
  .I1(sdpb_inst_115_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1538 (
  .O(mux_o_1538),
  .I0(sdpb_inst_116_dout[24]),
  .I1(sdpb_inst_117_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1539 (
  .O(mux_o_1539),
  .I0(sdpb_inst_118_dout[24]),
  .I1(sdpb_inst_119_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1540 (
  .O(mux_o_1540),
  .I0(sdpb_inst_120_dout[24]),
  .I1(sdpb_inst_121_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1541 (
  .O(mux_o_1541),
  .I0(sdpb_inst_122_dout[24]),
  .I1(sdpb_inst_123_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1542 (
  .O(mux_o_1542),
  .I0(sdpb_inst_124_dout[24]),
  .I1(sdpb_inst_125_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1543 (
  .O(mux_o_1543),
  .I0(sdpb_inst_126_dout[24]),
  .I1(sdpb_inst_127_dout[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1544 (
  .O(mux_o_1544),
  .I0(mux_o_1512),
  .I1(mux_o_1513),
  .S0(dff_q_4)
);
MUX2 mux_inst_1545 (
  .O(mux_o_1545),
  .I0(mux_o_1514),
  .I1(mux_o_1515),
  .S0(dff_q_4)
);
MUX2 mux_inst_1546 (
  .O(mux_o_1546),
  .I0(mux_o_1516),
  .I1(mux_o_1517),
  .S0(dff_q_4)
);
MUX2 mux_inst_1547 (
  .O(mux_o_1547),
  .I0(mux_o_1518),
  .I1(mux_o_1519),
  .S0(dff_q_4)
);
MUX2 mux_inst_1548 (
  .O(mux_o_1548),
  .I0(mux_o_1520),
  .I1(mux_o_1521),
  .S0(dff_q_4)
);
MUX2 mux_inst_1549 (
  .O(mux_o_1549),
  .I0(mux_o_1522),
  .I1(mux_o_1523),
  .S0(dff_q_4)
);
MUX2 mux_inst_1550 (
  .O(mux_o_1550),
  .I0(mux_o_1524),
  .I1(mux_o_1525),
  .S0(dff_q_4)
);
MUX2 mux_inst_1551 (
  .O(mux_o_1551),
  .I0(mux_o_1526),
  .I1(mux_o_1527),
  .S0(dff_q_4)
);
MUX2 mux_inst_1552 (
  .O(mux_o_1552),
  .I0(mux_o_1528),
  .I1(mux_o_1529),
  .S0(dff_q_4)
);
MUX2 mux_inst_1553 (
  .O(mux_o_1553),
  .I0(mux_o_1530),
  .I1(mux_o_1531),
  .S0(dff_q_4)
);
MUX2 mux_inst_1554 (
  .O(mux_o_1554),
  .I0(mux_o_1532),
  .I1(mux_o_1533),
  .S0(dff_q_4)
);
MUX2 mux_inst_1555 (
  .O(mux_o_1555),
  .I0(mux_o_1534),
  .I1(mux_o_1535),
  .S0(dff_q_4)
);
MUX2 mux_inst_1556 (
  .O(mux_o_1556),
  .I0(mux_o_1536),
  .I1(mux_o_1537),
  .S0(dff_q_4)
);
MUX2 mux_inst_1557 (
  .O(mux_o_1557),
  .I0(mux_o_1538),
  .I1(mux_o_1539),
  .S0(dff_q_4)
);
MUX2 mux_inst_1558 (
  .O(mux_o_1558),
  .I0(mux_o_1540),
  .I1(mux_o_1541),
  .S0(dff_q_4)
);
MUX2 mux_inst_1559 (
  .O(mux_o_1559),
  .I0(mux_o_1542),
  .I1(mux_o_1543),
  .S0(dff_q_4)
);
MUX2 mux_inst_1560 (
  .O(mux_o_1560),
  .I0(mux_o_1544),
  .I1(mux_o_1545),
  .S0(dff_q_3)
);
MUX2 mux_inst_1561 (
  .O(mux_o_1561),
  .I0(mux_o_1546),
  .I1(mux_o_1547),
  .S0(dff_q_3)
);
MUX2 mux_inst_1562 (
  .O(mux_o_1562),
  .I0(mux_o_1548),
  .I1(mux_o_1549),
  .S0(dff_q_3)
);
MUX2 mux_inst_1563 (
  .O(mux_o_1563),
  .I0(mux_o_1550),
  .I1(mux_o_1551),
  .S0(dff_q_3)
);
MUX2 mux_inst_1564 (
  .O(mux_o_1564),
  .I0(mux_o_1552),
  .I1(mux_o_1553),
  .S0(dff_q_3)
);
MUX2 mux_inst_1565 (
  .O(mux_o_1565),
  .I0(mux_o_1554),
  .I1(mux_o_1555),
  .S0(dff_q_3)
);
MUX2 mux_inst_1566 (
  .O(mux_o_1566),
  .I0(mux_o_1556),
  .I1(mux_o_1557),
  .S0(dff_q_3)
);
MUX2 mux_inst_1567 (
  .O(mux_o_1567),
  .I0(mux_o_1558),
  .I1(mux_o_1559),
  .S0(dff_q_3)
);
MUX2 mux_inst_1568 (
  .O(mux_o_1568),
  .I0(mux_o_1560),
  .I1(mux_o_1561),
  .S0(dff_q_2)
);
MUX2 mux_inst_1569 (
  .O(mux_o_1569),
  .I0(mux_o_1562),
  .I1(mux_o_1563),
  .S0(dff_q_2)
);
MUX2 mux_inst_1570 (
  .O(mux_o_1570),
  .I0(mux_o_1564),
  .I1(mux_o_1565),
  .S0(dff_q_2)
);
MUX2 mux_inst_1571 (
  .O(mux_o_1571),
  .I0(mux_o_1566),
  .I1(mux_o_1567),
  .S0(dff_q_2)
);
MUX2 mux_inst_1572 (
  .O(mux_o_1572),
  .I0(mux_o_1568),
  .I1(mux_o_1569),
  .S0(dff_q_1)
);
MUX2 mux_inst_1573 (
  .O(mux_o_1573),
  .I0(mux_o_1570),
  .I1(mux_o_1571),
  .S0(dff_q_1)
);
MUX2 mux_inst_1574 (
  .O(dout[24]),
  .I0(mux_o_1572),
  .I1(mux_o_1573),
  .S0(dff_q_0)
);
MUX2 mux_inst_1575 (
  .O(mux_o_1575),
  .I0(sdpb_inst_64_dout[25]),
  .I1(sdpb_inst_65_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1576 (
  .O(mux_o_1576),
  .I0(sdpb_inst_66_dout[25]),
  .I1(sdpb_inst_67_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1577 (
  .O(mux_o_1577),
  .I0(sdpb_inst_68_dout[25]),
  .I1(sdpb_inst_69_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1578 (
  .O(mux_o_1578),
  .I0(sdpb_inst_70_dout[25]),
  .I1(sdpb_inst_71_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1579 (
  .O(mux_o_1579),
  .I0(sdpb_inst_72_dout[25]),
  .I1(sdpb_inst_73_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1580 (
  .O(mux_o_1580),
  .I0(sdpb_inst_74_dout[25]),
  .I1(sdpb_inst_75_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1581 (
  .O(mux_o_1581),
  .I0(sdpb_inst_76_dout[25]),
  .I1(sdpb_inst_77_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1582 (
  .O(mux_o_1582),
  .I0(sdpb_inst_78_dout[25]),
  .I1(sdpb_inst_79_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1583 (
  .O(mux_o_1583),
  .I0(sdpb_inst_80_dout[25]),
  .I1(sdpb_inst_81_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1584 (
  .O(mux_o_1584),
  .I0(sdpb_inst_82_dout[25]),
  .I1(sdpb_inst_83_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1585 (
  .O(mux_o_1585),
  .I0(sdpb_inst_84_dout[25]),
  .I1(sdpb_inst_85_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1586 (
  .O(mux_o_1586),
  .I0(sdpb_inst_86_dout[25]),
  .I1(sdpb_inst_87_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1587 (
  .O(mux_o_1587),
  .I0(sdpb_inst_88_dout[25]),
  .I1(sdpb_inst_89_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1588 (
  .O(mux_o_1588),
  .I0(sdpb_inst_90_dout[25]),
  .I1(sdpb_inst_91_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1589 (
  .O(mux_o_1589),
  .I0(sdpb_inst_92_dout[25]),
  .I1(sdpb_inst_93_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1590 (
  .O(mux_o_1590),
  .I0(sdpb_inst_94_dout[25]),
  .I1(sdpb_inst_95_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1591 (
  .O(mux_o_1591),
  .I0(sdpb_inst_96_dout[25]),
  .I1(sdpb_inst_97_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1592 (
  .O(mux_o_1592),
  .I0(sdpb_inst_98_dout[25]),
  .I1(sdpb_inst_99_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1593 (
  .O(mux_o_1593),
  .I0(sdpb_inst_100_dout[25]),
  .I1(sdpb_inst_101_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1594 (
  .O(mux_o_1594),
  .I0(sdpb_inst_102_dout[25]),
  .I1(sdpb_inst_103_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1595 (
  .O(mux_o_1595),
  .I0(sdpb_inst_104_dout[25]),
  .I1(sdpb_inst_105_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1596 (
  .O(mux_o_1596),
  .I0(sdpb_inst_106_dout[25]),
  .I1(sdpb_inst_107_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1597 (
  .O(mux_o_1597),
  .I0(sdpb_inst_108_dout[25]),
  .I1(sdpb_inst_109_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1598 (
  .O(mux_o_1598),
  .I0(sdpb_inst_110_dout[25]),
  .I1(sdpb_inst_111_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1599 (
  .O(mux_o_1599),
  .I0(sdpb_inst_112_dout[25]),
  .I1(sdpb_inst_113_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1600 (
  .O(mux_o_1600),
  .I0(sdpb_inst_114_dout[25]),
  .I1(sdpb_inst_115_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1601 (
  .O(mux_o_1601),
  .I0(sdpb_inst_116_dout[25]),
  .I1(sdpb_inst_117_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1602 (
  .O(mux_o_1602),
  .I0(sdpb_inst_118_dout[25]),
  .I1(sdpb_inst_119_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1603 (
  .O(mux_o_1603),
  .I0(sdpb_inst_120_dout[25]),
  .I1(sdpb_inst_121_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1604 (
  .O(mux_o_1604),
  .I0(sdpb_inst_122_dout[25]),
  .I1(sdpb_inst_123_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1605 (
  .O(mux_o_1605),
  .I0(sdpb_inst_124_dout[25]),
  .I1(sdpb_inst_125_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1606 (
  .O(mux_o_1606),
  .I0(sdpb_inst_126_dout[25]),
  .I1(sdpb_inst_127_dout[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1607 (
  .O(mux_o_1607),
  .I0(mux_o_1575),
  .I1(mux_o_1576),
  .S0(dff_q_4)
);
MUX2 mux_inst_1608 (
  .O(mux_o_1608),
  .I0(mux_o_1577),
  .I1(mux_o_1578),
  .S0(dff_q_4)
);
MUX2 mux_inst_1609 (
  .O(mux_o_1609),
  .I0(mux_o_1579),
  .I1(mux_o_1580),
  .S0(dff_q_4)
);
MUX2 mux_inst_1610 (
  .O(mux_o_1610),
  .I0(mux_o_1581),
  .I1(mux_o_1582),
  .S0(dff_q_4)
);
MUX2 mux_inst_1611 (
  .O(mux_o_1611),
  .I0(mux_o_1583),
  .I1(mux_o_1584),
  .S0(dff_q_4)
);
MUX2 mux_inst_1612 (
  .O(mux_o_1612),
  .I0(mux_o_1585),
  .I1(mux_o_1586),
  .S0(dff_q_4)
);
MUX2 mux_inst_1613 (
  .O(mux_o_1613),
  .I0(mux_o_1587),
  .I1(mux_o_1588),
  .S0(dff_q_4)
);
MUX2 mux_inst_1614 (
  .O(mux_o_1614),
  .I0(mux_o_1589),
  .I1(mux_o_1590),
  .S0(dff_q_4)
);
MUX2 mux_inst_1615 (
  .O(mux_o_1615),
  .I0(mux_o_1591),
  .I1(mux_o_1592),
  .S0(dff_q_4)
);
MUX2 mux_inst_1616 (
  .O(mux_o_1616),
  .I0(mux_o_1593),
  .I1(mux_o_1594),
  .S0(dff_q_4)
);
MUX2 mux_inst_1617 (
  .O(mux_o_1617),
  .I0(mux_o_1595),
  .I1(mux_o_1596),
  .S0(dff_q_4)
);
MUX2 mux_inst_1618 (
  .O(mux_o_1618),
  .I0(mux_o_1597),
  .I1(mux_o_1598),
  .S0(dff_q_4)
);
MUX2 mux_inst_1619 (
  .O(mux_o_1619),
  .I0(mux_o_1599),
  .I1(mux_o_1600),
  .S0(dff_q_4)
);
MUX2 mux_inst_1620 (
  .O(mux_o_1620),
  .I0(mux_o_1601),
  .I1(mux_o_1602),
  .S0(dff_q_4)
);
MUX2 mux_inst_1621 (
  .O(mux_o_1621),
  .I0(mux_o_1603),
  .I1(mux_o_1604),
  .S0(dff_q_4)
);
MUX2 mux_inst_1622 (
  .O(mux_o_1622),
  .I0(mux_o_1605),
  .I1(mux_o_1606),
  .S0(dff_q_4)
);
MUX2 mux_inst_1623 (
  .O(mux_o_1623),
  .I0(mux_o_1607),
  .I1(mux_o_1608),
  .S0(dff_q_3)
);
MUX2 mux_inst_1624 (
  .O(mux_o_1624),
  .I0(mux_o_1609),
  .I1(mux_o_1610),
  .S0(dff_q_3)
);
MUX2 mux_inst_1625 (
  .O(mux_o_1625),
  .I0(mux_o_1611),
  .I1(mux_o_1612),
  .S0(dff_q_3)
);
MUX2 mux_inst_1626 (
  .O(mux_o_1626),
  .I0(mux_o_1613),
  .I1(mux_o_1614),
  .S0(dff_q_3)
);
MUX2 mux_inst_1627 (
  .O(mux_o_1627),
  .I0(mux_o_1615),
  .I1(mux_o_1616),
  .S0(dff_q_3)
);
MUX2 mux_inst_1628 (
  .O(mux_o_1628),
  .I0(mux_o_1617),
  .I1(mux_o_1618),
  .S0(dff_q_3)
);
MUX2 mux_inst_1629 (
  .O(mux_o_1629),
  .I0(mux_o_1619),
  .I1(mux_o_1620),
  .S0(dff_q_3)
);
MUX2 mux_inst_1630 (
  .O(mux_o_1630),
  .I0(mux_o_1621),
  .I1(mux_o_1622),
  .S0(dff_q_3)
);
MUX2 mux_inst_1631 (
  .O(mux_o_1631),
  .I0(mux_o_1623),
  .I1(mux_o_1624),
  .S0(dff_q_2)
);
MUX2 mux_inst_1632 (
  .O(mux_o_1632),
  .I0(mux_o_1625),
  .I1(mux_o_1626),
  .S0(dff_q_2)
);
MUX2 mux_inst_1633 (
  .O(mux_o_1633),
  .I0(mux_o_1627),
  .I1(mux_o_1628),
  .S0(dff_q_2)
);
MUX2 mux_inst_1634 (
  .O(mux_o_1634),
  .I0(mux_o_1629),
  .I1(mux_o_1630),
  .S0(dff_q_2)
);
MUX2 mux_inst_1635 (
  .O(mux_o_1635),
  .I0(mux_o_1631),
  .I1(mux_o_1632),
  .S0(dff_q_1)
);
MUX2 mux_inst_1636 (
  .O(mux_o_1636),
  .I0(mux_o_1633),
  .I1(mux_o_1634),
  .S0(dff_q_1)
);
MUX2 mux_inst_1637 (
  .O(dout[25]),
  .I0(mux_o_1635),
  .I1(mux_o_1636),
  .S0(dff_q_0)
);
MUX2 mux_inst_1638 (
  .O(mux_o_1638),
  .I0(sdpb_inst_64_dout[26]),
  .I1(sdpb_inst_65_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1639 (
  .O(mux_o_1639),
  .I0(sdpb_inst_66_dout[26]),
  .I1(sdpb_inst_67_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1640 (
  .O(mux_o_1640),
  .I0(sdpb_inst_68_dout[26]),
  .I1(sdpb_inst_69_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1641 (
  .O(mux_o_1641),
  .I0(sdpb_inst_70_dout[26]),
  .I1(sdpb_inst_71_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1642 (
  .O(mux_o_1642),
  .I0(sdpb_inst_72_dout[26]),
  .I1(sdpb_inst_73_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1643 (
  .O(mux_o_1643),
  .I0(sdpb_inst_74_dout[26]),
  .I1(sdpb_inst_75_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1644 (
  .O(mux_o_1644),
  .I0(sdpb_inst_76_dout[26]),
  .I1(sdpb_inst_77_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1645 (
  .O(mux_o_1645),
  .I0(sdpb_inst_78_dout[26]),
  .I1(sdpb_inst_79_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1646 (
  .O(mux_o_1646),
  .I0(sdpb_inst_80_dout[26]),
  .I1(sdpb_inst_81_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1647 (
  .O(mux_o_1647),
  .I0(sdpb_inst_82_dout[26]),
  .I1(sdpb_inst_83_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1648 (
  .O(mux_o_1648),
  .I0(sdpb_inst_84_dout[26]),
  .I1(sdpb_inst_85_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1649 (
  .O(mux_o_1649),
  .I0(sdpb_inst_86_dout[26]),
  .I1(sdpb_inst_87_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1650 (
  .O(mux_o_1650),
  .I0(sdpb_inst_88_dout[26]),
  .I1(sdpb_inst_89_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1651 (
  .O(mux_o_1651),
  .I0(sdpb_inst_90_dout[26]),
  .I1(sdpb_inst_91_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1652 (
  .O(mux_o_1652),
  .I0(sdpb_inst_92_dout[26]),
  .I1(sdpb_inst_93_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1653 (
  .O(mux_o_1653),
  .I0(sdpb_inst_94_dout[26]),
  .I1(sdpb_inst_95_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1654 (
  .O(mux_o_1654),
  .I0(sdpb_inst_96_dout[26]),
  .I1(sdpb_inst_97_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1655 (
  .O(mux_o_1655),
  .I0(sdpb_inst_98_dout[26]),
  .I1(sdpb_inst_99_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1656 (
  .O(mux_o_1656),
  .I0(sdpb_inst_100_dout[26]),
  .I1(sdpb_inst_101_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1657 (
  .O(mux_o_1657),
  .I0(sdpb_inst_102_dout[26]),
  .I1(sdpb_inst_103_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1658 (
  .O(mux_o_1658),
  .I0(sdpb_inst_104_dout[26]),
  .I1(sdpb_inst_105_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1659 (
  .O(mux_o_1659),
  .I0(sdpb_inst_106_dout[26]),
  .I1(sdpb_inst_107_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1660 (
  .O(mux_o_1660),
  .I0(sdpb_inst_108_dout[26]),
  .I1(sdpb_inst_109_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1661 (
  .O(mux_o_1661),
  .I0(sdpb_inst_110_dout[26]),
  .I1(sdpb_inst_111_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1662 (
  .O(mux_o_1662),
  .I0(sdpb_inst_112_dout[26]),
  .I1(sdpb_inst_113_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1663 (
  .O(mux_o_1663),
  .I0(sdpb_inst_114_dout[26]),
  .I1(sdpb_inst_115_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1664 (
  .O(mux_o_1664),
  .I0(sdpb_inst_116_dout[26]),
  .I1(sdpb_inst_117_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1665 (
  .O(mux_o_1665),
  .I0(sdpb_inst_118_dout[26]),
  .I1(sdpb_inst_119_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1666 (
  .O(mux_o_1666),
  .I0(sdpb_inst_120_dout[26]),
  .I1(sdpb_inst_121_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1667 (
  .O(mux_o_1667),
  .I0(sdpb_inst_122_dout[26]),
  .I1(sdpb_inst_123_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1668 (
  .O(mux_o_1668),
  .I0(sdpb_inst_124_dout[26]),
  .I1(sdpb_inst_125_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1669 (
  .O(mux_o_1669),
  .I0(sdpb_inst_126_dout[26]),
  .I1(sdpb_inst_127_dout[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1670 (
  .O(mux_o_1670),
  .I0(mux_o_1638),
  .I1(mux_o_1639),
  .S0(dff_q_4)
);
MUX2 mux_inst_1671 (
  .O(mux_o_1671),
  .I0(mux_o_1640),
  .I1(mux_o_1641),
  .S0(dff_q_4)
);
MUX2 mux_inst_1672 (
  .O(mux_o_1672),
  .I0(mux_o_1642),
  .I1(mux_o_1643),
  .S0(dff_q_4)
);
MUX2 mux_inst_1673 (
  .O(mux_o_1673),
  .I0(mux_o_1644),
  .I1(mux_o_1645),
  .S0(dff_q_4)
);
MUX2 mux_inst_1674 (
  .O(mux_o_1674),
  .I0(mux_o_1646),
  .I1(mux_o_1647),
  .S0(dff_q_4)
);
MUX2 mux_inst_1675 (
  .O(mux_o_1675),
  .I0(mux_o_1648),
  .I1(mux_o_1649),
  .S0(dff_q_4)
);
MUX2 mux_inst_1676 (
  .O(mux_o_1676),
  .I0(mux_o_1650),
  .I1(mux_o_1651),
  .S0(dff_q_4)
);
MUX2 mux_inst_1677 (
  .O(mux_o_1677),
  .I0(mux_o_1652),
  .I1(mux_o_1653),
  .S0(dff_q_4)
);
MUX2 mux_inst_1678 (
  .O(mux_o_1678),
  .I0(mux_o_1654),
  .I1(mux_o_1655),
  .S0(dff_q_4)
);
MUX2 mux_inst_1679 (
  .O(mux_o_1679),
  .I0(mux_o_1656),
  .I1(mux_o_1657),
  .S0(dff_q_4)
);
MUX2 mux_inst_1680 (
  .O(mux_o_1680),
  .I0(mux_o_1658),
  .I1(mux_o_1659),
  .S0(dff_q_4)
);
MUX2 mux_inst_1681 (
  .O(mux_o_1681),
  .I0(mux_o_1660),
  .I1(mux_o_1661),
  .S0(dff_q_4)
);
MUX2 mux_inst_1682 (
  .O(mux_o_1682),
  .I0(mux_o_1662),
  .I1(mux_o_1663),
  .S0(dff_q_4)
);
MUX2 mux_inst_1683 (
  .O(mux_o_1683),
  .I0(mux_o_1664),
  .I1(mux_o_1665),
  .S0(dff_q_4)
);
MUX2 mux_inst_1684 (
  .O(mux_o_1684),
  .I0(mux_o_1666),
  .I1(mux_o_1667),
  .S0(dff_q_4)
);
MUX2 mux_inst_1685 (
  .O(mux_o_1685),
  .I0(mux_o_1668),
  .I1(mux_o_1669),
  .S0(dff_q_4)
);
MUX2 mux_inst_1686 (
  .O(mux_o_1686),
  .I0(mux_o_1670),
  .I1(mux_o_1671),
  .S0(dff_q_3)
);
MUX2 mux_inst_1687 (
  .O(mux_o_1687),
  .I0(mux_o_1672),
  .I1(mux_o_1673),
  .S0(dff_q_3)
);
MUX2 mux_inst_1688 (
  .O(mux_o_1688),
  .I0(mux_o_1674),
  .I1(mux_o_1675),
  .S0(dff_q_3)
);
MUX2 mux_inst_1689 (
  .O(mux_o_1689),
  .I0(mux_o_1676),
  .I1(mux_o_1677),
  .S0(dff_q_3)
);
MUX2 mux_inst_1690 (
  .O(mux_o_1690),
  .I0(mux_o_1678),
  .I1(mux_o_1679),
  .S0(dff_q_3)
);
MUX2 mux_inst_1691 (
  .O(mux_o_1691),
  .I0(mux_o_1680),
  .I1(mux_o_1681),
  .S0(dff_q_3)
);
MUX2 mux_inst_1692 (
  .O(mux_o_1692),
  .I0(mux_o_1682),
  .I1(mux_o_1683),
  .S0(dff_q_3)
);
MUX2 mux_inst_1693 (
  .O(mux_o_1693),
  .I0(mux_o_1684),
  .I1(mux_o_1685),
  .S0(dff_q_3)
);
MUX2 mux_inst_1694 (
  .O(mux_o_1694),
  .I0(mux_o_1686),
  .I1(mux_o_1687),
  .S0(dff_q_2)
);
MUX2 mux_inst_1695 (
  .O(mux_o_1695),
  .I0(mux_o_1688),
  .I1(mux_o_1689),
  .S0(dff_q_2)
);
MUX2 mux_inst_1696 (
  .O(mux_o_1696),
  .I0(mux_o_1690),
  .I1(mux_o_1691),
  .S0(dff_q_2)
);
MUX2 mux_inst_1697 (
  .O(mux_o_1697),
  .I0(mux_o_1692),
  .I1(mux_o_1693),
  .S0(dff_q_2)
);
MUX2 mux_inst_1698 (
  .O(mux_o_1698),
  .I0(mux_o_1694),
  .I1(mux_o_1695),
  .S0(dff_q_1)
);
MUX2 mux_inst_1699 (
  .O(mux_o_1699),
  .I0(mux_o_1696),
  .I1(mux_o_1697),
  .S0(dff_q_1)
);
MUX2 mux_inst_1700 (
  .O(dout[26]),
  .I0(mux_o_1698),
  .I1(mux_o_1699),
  .S0(dff_q_0)
);
MUX2 mux_inst_1701 (
  .O(mux_o_1701),
  .I0(sdpb_inst_64_dout[27]),
  .I1(sdpb_inst_65_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1702 (
  .O(mux_o_1702),
  .I0(sdpb_inst_66_dout[27]),
  .I1(sdpb_inst_67_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1703 (
  .O(mux_o_1703),
  .I0(sdpb_inst_68_dout[27]),
  .I1(sdpb_inst_69_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1704 (
  .O(mux_o_1704),
  .I0(sdpb_inst_70_dout[27]),
  .I1(sdpb_inst_71_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1705 (
  .O(mux_o_1705),
  .I0(sdpb_inst_72_dout[27]),
  .I1(sdpb_inst_73_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1706 (
  .O(mux_o_1706),
  .I0(sdpb_inst_74_dout[27]),
  .I1(sdpb_inst_75_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1707 (
  .O(mux_o_1707),
  .I0(sdpb_inst_76_dout[27]),
  .I1(sdpb_inst_77_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1708 (
  .O(mux_o_1708),
  .I0(sdpb_inst_78_dout[27]),
  .I1(sdpb_inst_79_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1709 (
  .O(mux_o_1709),
  .I0(sdpb_inst_80_dout[27]),
  .I1(sdpb_inst_81_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1710 (
  .O(mux_o_1710),
  .I0(sdpb_inst_82_dout[27]),
  .I1(sdpb_inst_83_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1711 (
  .O(mux_o_1711),
  .I0(sdpb_inst_84_dout[27]),
  .I1(sdpb_inst_85_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1712 (
  .O(mux_o_1712),
  .I0(sdpb_inst_86_dout[27]),
  .I1(sdpb_inst_87_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1713 (
  .O(mux_o_1713),
  .I0(sdpb_inst_88_dout[27]),
  .I1(sdpb_inst_89_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1714 (
  .O(mux_o_1714),
  .I0(sdpb_inst_90_dout[27]),
  .I1(sdpb_inst_91_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1715 (
  .O(mux_o_1715),
  .I0(sdpb_inst_92_dout[27]),
  .I1(sdpb_inst_93_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1716 (
  .O(mux_o_1716),
  .I0(sdpb_inst_94_dout[27]),
  .I1(sdpb_inst_95_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1717 (
  .O(mux_o_1717),
  .I0(sdpb_inst_96_dout[27]),
  .I1(sdpb_inst_97_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1718 (
  .O(mux_o_1718),
  .I0(sdpb_inst_98_dout[27]),
  .I1(sdpb_inst_99_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1719 (
  .O(mux_o_1719),
  .I0(sdpb_inst_100_dout[27]),
  .I1(sdpb_inst_101_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1720 (
  .O(mux_o_1720),
  .I0(sdpb_inst_102_dout[27]),
  .I1(sdpb_inst_103_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1721 (
  .O(mux_o_1721),
  .I0(sdpb_inst_104_dout[27]),
  .I1(sdpb_inst_105_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1722 (
  .O(mux_o_1722),
  .I0(sdpb_inst_106_dout[27]),
  .I1(sdpb_inst_107_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1723 (
  .O(mux_o_1723),
  .I0(sdpb_inst_108_dout[27]),
  .I1(sdpb_inst_109_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1724 (
  .O(mux_o_1724),
  .I0(sdpb_inst_110_dout[27]),
  .I1(sdpb_inst_111_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1725 (
  .O(mux_o_1725),
  .I0(sdpb_inst_112_dout[27]),
  .I1(sdpb_inst_113_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1726 (
  .O(mux_o_1726),
  .I0(sdpb_inst_114_dout[27]),
  .I1(sdpb_inst_115_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1727 (
  .O(mux_o_1727),
  .I0(sdpb_inst_116_dout[27]),
  .I1(sdpb_inst_117_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1728 (
  .O(mux_o_1728),
  .I0(sdpb_inst_118_dout[27]),
  .I1(sdpb_inst_119_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1729 (
  .O(mux_o_1729),
  .I0(sdpb_inst_120_dout[27]),
  .I1(sdpb_inst_121_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1730 (
  .O(mux_o_1730),
  .I0(sdpb_inst_122_dout[27]),
  .I1(sdpb_inst_123_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1731 (
  .O(mux_o_1731),
  .I0(sdpb_inst_124_dout[27]),
  .I1(sdpb_inst_125_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1732 (
  .O(mux_o_1732),
  .I0(sdpb_inst_126_dout[27]),
  .I1(sdpb_inst_127_dout[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1733 (
  .O(mux_o_1733),
  .I0(mux_o_1701),
  .I1(mux_o_1702),
  .S0(dff_q_4)
);
MUX2 mux_inst_1734 (
  .O(mux_o_1734),
  .I0(mux_o_1703),
  .I1(mux_o_1704),
  .S0(dff_q_4)
);
MUX2 mux_inst_1735 (
  .O(mux_o_1735),
  .I0(mux_o_1705),
  .I1(mux_o_1706),
  .S0(dff_q_4)
);
MUX2 mux_inst_1736 (
  .O(mux_o_1736),
  .I0(mux_o_1707),
  .I1(mux_o_1708),
  .S0(dff_q_4)
);
MUX2 mux_inst_1737 (
  .O(mux_o_1737),
  .I0(mux_o_1709),
  .I1(mux_o_1710),
  .S0(dff_q_4)
);
MUX2 mux_inst_1738 (
  .O(mux_o_1738),
  .I0(mux_o_1711),
  .I1(mux_o_1712),
  .S0(dff_q_4)
);
MUX2 mux_inst_1739 (
  .O(mux_o_1739),
  .I0(mux_o_1713),
  .I1(mux_o_1714),
  .S0(dff_q_4)
);
MUX2 mux_inst_1740 (
  .O(mux_o_1740),
  .I0(mux_o_1715),
  .I1(mux_o_1716),
  .S0(dff_q_4)
);
MUX2 mux_inst_1741 (
  .O(mux_o_1741),
  .I0(mux_o_1717),
  .I1(mux_o_1718),
  .S0(dff_q_4)
);
MUX2 mux_inst_1742 (
  .O(mux_o_1742),
  .I0(mux_o_1719),
  .I1(mux_o_1720),
  .S0(dff_q_4)
);
MUX2 mux_inst_1743 (
  .O(mux_o_1743),
  .I0(mux_o_1721),
  .I1(mux_o_1722),
  .S0(dff_q_4)
);
MUX2 mux_inst_1744 (
  .O(mux_o_1744),
  .I0(mux_o_1723),
  .I1(mux_o_1724),
  .S0(dff_q_4)
);
MUX2 mux_inst_1745 (
  .O(mux_o_1745),
  .I0(mux_o_1725),
  .I1(mux_o_1726),
  .S0(dff_q_4)
);
MUX2 mux_inst_1746 (
  .O(mux_o_1746),
  .I0(mux_o_1727),
  .I1(mux_o_1728),
  .S0(dff_q_4)
);
MUX2 mux_inst_1747 (
  .O(mux_o_1747),
  .I0(mux_o_1729),
  .I1(mux_o_1730),
  .S0(dff_q_4)
);
MUX2 mux_inst_1748 (
  .O(mux_o_1748),
  .I0(mux_o_1731),
  .I1(mux_o_1732),
  .S0(dff_q_4)
);
MUX2 mux_inst_1749 (
  .O(mux_o_1749),
  .I0(mux_o_1733),
  .I1(mux_o_1734),
  .S0(dff_q_3)
);
MUX2 mux_inst_1750 (
  .O(mux_o_1750),
  .I0(mux_o_1735),
  .I1(mux_o_1736),
  .S0(dff_q_3)
);
MUX2 mux_inst_1751 (
  .O(mux_o_1751),
  .I0(mux_o_1737),
  .I1(mux_o_1738),
  .S0(dff_q_3)
);
MUX2 mux_inst_1752 (
  .O(mux_o_1752),
  .I0(mux_o_1739),
  .I1(mux_o_1740),
  .S0(dff_q_3)
);
MUX2 mux_inst_1753 (
  .O(mux_o_1753),
  .I0(mux_o_1741),
  .I1(mux_o_1742),
  .S0(dff_q_3)
);
MUX2 mux_inst_1754 (
  .O(mux_o_1754),
  .I0(mux_o_1743),
  .I1(mux_o_1744),
  .S0(dff_q_3)
);
MUX2 mux_inst_1755 (
  .O(mux_o_1755),
  .I0(mux_o_1745),
  .I1(mux_o_1746),
  .S0(dff_q_3)
);
MUX2 mux_inst_1756 (
  .O(mux_o_1756),
  .I0(mux_o_1747),
  .I1(mux_o_1748),
  .S0(dff_q_3)
);
MUX2 mux_inst_1757 (
  .O(mux_o_1757),
  .I0(mux_o_1749),
  .I1(mux_o_1750),
  .S0(dff_q_2)
);
MUX2 mux_inst_1758 (
  .O(mux_o_1758),
  .I0(mux_o_1751),
  .I1(mux_o_1752),
  .S0(dff_q_2)
);
MUX2 mux_inst_1759 (
  .O(mux_o_1759),
  .I0(mux_o_1753),
  .I1(mux_o_1754),
  .S0(dff_q_2)
);
MUX2 mux_inst_1760 (
  .O(mux_o_1760),
  .I0(mux_o_1755),
  .I1(mux_o_1756),
  .S0(dff_q_2)
);
MUX2 mux_inst_1761 (
  .O(mux_o_1761),
  .I0(mux_o_1757),
  .I1(mux_o_1758),
  .S0(dff_q_1)
);
MUX2 mux_inst_1762 (
  .O(mux_o_1762),
  .I0(mux_o_1759),
  .I1(mux_o_1760),
  .S0(dff_q_1)
);
MUX2 mux_inst_1763 (
  .O(dout[27]),
  .I0(mux_o_1761),
  .I1(mux_o_1762),
  .S0(dff_q_0)
);
MUX2 mux_inst_1764 (
  .O(mux_o_1764),
  .I0(sdpb_inst_64_dout[28]),
  .I1(sdpb_inst_65_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1765 (
  .O(mux_o_1765),
  .I0(sdpb_inst_66_dout[28]),
  .I1(sdpb_inst_67_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1766 (
  .O(mux_o_1766),
  .I0(sdpb_inst_68_dout[28]),
  .I1(sdpb_inst_69_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1767 (
  .O(mux_o_1767),
  .I0(sdpb_inst_70_dout[28]),
  .I1(sdpb_inst_71_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1768 (
  .O(mux_o_1768),
  .I0(sdpb_inst_72_dout[28]),
  .I1(sdpb_inst_73_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1769 (
  .O(mux_o_1769),
  .I0(sdpb_inst_74_dout[28]),
  .I1(sdpb_inst_75_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1770 (
  .O(mux_o_1770),
  .I0(sdpb_inst_76_dout[28]),
  .I1(sdpb_inst_77_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1771 (
  .O(mux_o_1771),
  .I0(sdpb_inst_78_dout[28]),
  .I1(sdpb_inst_79_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1772 (
  .O(mux_o_1772),
  .I0(sdpb_inst_80_dout[28]),
  .I1(sdpb_inst_81_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1773 (
  .O(mux_o_1773),
  .I0(sdpb_inst_82_dout[28]),
  .I1(sdpb_inst_83_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1774 (
  .O(mux_o_1774),
  .I0(sdpb_inst_84_dout[28]),
  .I1(sdpb_inst_85_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1775 (
  .O(mux_o_1775),
  .I0(sdpb_inst_86_dout[28]),
  .I1(sdpb_inst_87_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1776 (
  .O(mux_o_1776),
  .I0(sdpb_inst_88_dout[28]),
  .I1(sdpb_inst_89_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1777 (
  .O(mux_o_1777),
  .I0(sdpb_inst_90_dout[28]),
  .I1(sdpb_inst_91_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1778 (
  .O(mux_o_1778),
  .I0(sdpb_inst_92_dout[28]),
  .I1(sdpb_inst_93_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1779 (
  .O(mux_o_1779),
  .I0(sdpb_inst_94_dout[28]),
  .I1(sdpb_inst_95_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1780 (
  .O(mux_o_1780),
  .I0(sdpb_inst_96_dout[28]),
  .I1(sdpb_inst_97_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1781 (
  .O(mux_o_1781),
  .I0(sdpb_inst_98_dout[28]),
  .I1(sdpb_inst_99_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1782 (
  .O(mux_o_1782),
  .I0(sdpb_inst_100_dout[28]),
  .I1(sdpb_inst_101_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1783 (
  .O(mux_o_1783),
  .I0(sdpb_inst_102_dout[28]),
  .I1(sdpb_inst_103_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1784 (
  .O(mux_o_1784),
  .I0(sdpb_inst_104_dout[28]),
  .I1(sdpb_inst_105_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1785 (
  .O(mux_o_1785),
  .I0(sdpb_inst_106_dout[28]),
  .I1(sdpb_inst_107_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1786 (
  .O(mux_o_1786),
  .I0(sdpb_inst_108_dout[28]),
  .I1(sdpb_inst_109_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1787 (
  .O(mux_o_1787),
  .I0(sdpb_inst_110_dout[28]),
  .I1(sdpb_inst_111_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1788 (
  .O(mux_o_1788),
  .I0(sdpb_inst_112_dout[28]),
  .I1(sdpb_inst_113_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1789 (
  .O(mux_o_1789),
  .I0(sdpb_inst_114_dout[28]),
  .I1(sdpb_inst_115_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1790 (
  .O(mux_o_1790),
  .I0(sdpb_inst_116_dout[28]),
  .I1(sdpb_inst_117_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1791 (
  .O(mux_o_1791),
  .I0(sdpb_inst_118_dout[28]),
  .I1(sdpb_inst_119_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1792 (
  .O(mux_o_1792),
  .I0(sdpb_inst_120_dout[28]),
  .I1(sdpb_inst_121_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1793 (
  .O(mux_o_1793),
  .I0(sdpb_inst_122_dout[28]),
  .I1(sdpb_inst_123_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1794 (
  .O(mux_o_1794),
  .I0(sdpb_inst_124_dout[28]),
  .I1(sdpb_inst_125_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1795 (
  .O(mux_o_1795),
  .I0(sdpb_inst_126_dout[28]),
  .I1(sdpb_inst_127_dout[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1796 (
  .O(mux_o_1796),
  .I0(mux_o_1764),
  .I1(mux_o_1765),
  .S0(dff_q_4)
);
MUX2 mux_inst_1797 (
  .O(mux_o_1797),
  .I0(mux_o_1766),
  .I1(mux_o_1767),
  .S0(dff_q_4)
);
MUX2 mux_inst_1798 (
  .O(mux_o_1798),
  .I0(mux_o_1768),
  .I1(mux_o_1769),
  .S0(dff_q_4)
);
MUX2 mux_inst_1799 (
  .O(mux_o_1799),
  .I0(mux_o_1770),
  .I1(mux_o_1771),
  .S0(dff_q_4)
);
MUX2 mux_inst_1800 (
  .O(mux_o_1800),
  .I0(mux_o_1772),
  .I1(mux_o_1773),
  .S0(dff_q_4)
);
MUX2 mux_inst_1801 (
  .O(mux_o_1801),
  .I0(mux_o_1774),
  .I1(mux_o_1775),
  .S0(dff_q_4)
);
MUX2 mux_inst_1802 (
  .O(mux_o_1802),
  .I0(mux_o_1776),
  .I1(mux_o_1777),
  .S0(dff_q_4)
);
MUX2 mux_inst_1803 (
  .O(mux_o_1803),
  .I0(mux_o_1778),
  .I1(mux_o_1779),
  .S0(dff_q_4)
);
MUX2 mux_inst_1804 (
  .O(mux_o_1804),
  .I0(mux_o_1780),
  .I1(mux_o_1781),
  .S0(dff_q_4)
);
MUX2 mux_inst_1805 (
  .O(mux_o_1805),
  .I0(mux_o_1782),
  .I1(mux_o_1783),
  .S0(dff_q_4)
);
MUX2 mux_inst_1806 (
  .O(mux_o_1806),
  .I0(mux_o_1784),
  .I1(mux_o_1785),
  .S0(dff_q_4)
);
MUX2 mux_inst_1807 (
  .O(mux_o_1807),
  .I0(mux_o_1786),
  .I1(mux_o_1787),
  .S0(dff_q_4)
);
MUX2 mux_inst_1808 (
  .O(mux_o_1808),
  .I0(mux_o_1788),
  .I1(mux_o_1789),
  .S0(dff_q_4)
);
MUX2 mux_inst_1809 (
  .O(mux_o_1809),
  .I0(mux_o_1790),
  .I1(mux_o_1791),
  .S0(dff_q_4)
);
MUX2 mux_inst_1810 (
  .O(mux_o_1810),
  .I0(mux_o_1792),
  .I1(mux_o_1793),
  .S0(dff_q_4)
);
MUX2 mux_inst_1811 (
  .O(mux_o_1811),
  .I0(mux_o_1794),
  .I1(mux_o_1795),
  .S0(dff_q_4)
);
MUX2 mux_inst_1812 (
  .O(mux_o_1812),
  .I0(mux_o_1796),
  .I1(mux_o_1797),
  .S0(dff_q_3)
);
MUX2 mux_inst_1813 (
  .O(mux_o_1813),
  .I0(mux_o_1798),
  .I1(mux_o_1799),
  .S0(dff_q_3)
);
MUX2 mux_inst_1814 (
  .O(mux_o_1814),
  .I0(mux_o_1800),
  .I1(mux_o_1801),
  .S0(dff_q_3)
);
MUX2 mux_inst_1815 (
  .O(mux_o_1815),
  .I0(mux_o_1802),
  .I1(mux_o_1803),
  .S0(dff_q_3)
);
MUX2 mux_inst_1816 (
  .O(mux_o_1816),
  .I0(mux_o_1804),
  .I1(mux_o_1805),
  .S0(dff_q_3)
);
MUX2 mux_inst_1817 (
  .O(mux_o_1817),
  .I0(mux_o_1806),
  .I1(mux_o_1807),
  .S0(dff_q_3)
);
MUX2 mux_inst_1818 (
  .O(mux_o_1818),
  .I0(mux_o_1808),
  .I1(mux_o_1809),
  .S0(dff_q_3)
);
MUX2 mux_inst_1819 (
  .O(mux_o_1819),
  .I0(mux_o_1810),
  .I1(mux_o_1811),
  .S0(dff_q_3)
);
MUX2 mux_inst_1820 (
  .O(mux_o_1820),
  .I0(mux_o_1812),
  .I1(mux_o_1813),
  .S0(dff_q_2)
);
MUX2 mux_inst_1821 (
  .O(mux_o_1821),
  .I0(mux_o_1814),
  .I1(mux_o_1815),
  .S0(dff_q_2)
);
MUX2 mux_inst_1822 (
  .O(mux_o_1822),
  .I0(mux_o_1816),
  .I1(mux_o_1817),
  .S0(dff_q_2)
);
MUX2 mux_inst_1823 (
  .O(mux_o_1823),
  .I0(mux_o_1818),
  .I1(mux_o_1819),
  .S0(dff_q_2)
);
MUX2 mux_inst_1824 (
  .O(mux_o_1824),
  .I0(mux_o_1820),
  .I1(mux_o_1821),
  .S0(dff_q_1)
);
MUX2 mux_inst_1825 (
  .O(mux_o_1825),
  .I0(mux_o_1822),
  .I1(mux_o_1823),
  .S0(dff_q_1)
);
MUX2 mux_inst_1826 (
  .O(dout[28]),
  .I0(mux_o_1824),
  .I1(mux_o_1825),
  .S0(dff_q_0)
);
MUX2 mux_inst_1827 (
  .O(mux_o_1827),
  .I0(sdpb_inst_64_dout[29]),
  .I1(sdpb_inst_65_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1828 (
  .O(mux_o_1828),
  .I0(sdpb_inst_66_dout[29]),
  .I1(sdpb_inst_67_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1829 (
  .O(mux_o_1829),
  .I0(sdpb_inst_68_dout[29]),
  .I1(sdpb_inst_69_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1830 (
  .O(mux_o_1830),
  .I0(sdpb_inst_70_dout[29]),
  .I1(sdpb_inst_71_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1831 (
  .O(mux_o_1831),
  .I0(sdpb_inst_72_dout[29]),
  .I1(sdpb_inst_73_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1832 (
  .O(mux_o_1832),
  .I0(sdpb_inst_74_dout[29]),
  .I1(sdpb_inst_75_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1833 (
  .O(mux_o_1833),
  .I0(sdpb_inst_76_dout[29]),
  .I1(sdpb_inst_77_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1834 (
  .O(mux_o_1834),
  .I0(sdpb_inst_78_dout[29]),
  .I1(sdpb_inst_79_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1835 (
  .O(mux_o_1835),
  .I0(sdpb_inst_80_dout[29]),
  .I1(sdpb_inst_81_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1836 (
  .O(mux_o_1836),
  .I0(sdpb_inst_82_dout[29]),
  .I1(sdpb_inst_83_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1837 (
  .O(mux_o_1837),
  .I0(sdpb_inst_84_dout[29]),
  .I1(sdpb_inst_85_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1838 (
  .O(mux_o_1838),
  .I0(sdpb_inst_86_dout[29]),
  .I1(sdpb_inst_87_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1839 (
  .O(mux_o_1839),
  .I0(sdpb_inst_88_dout[29]),
  .I1(sdpb_inst_89_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1840 (
  .O(mux_o_1840),
  .I0(sdpb_inst_90_dout[29]),
  .I1(sdpb_inst_91_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1841 (
  .O(mux_o_1841),
  .I0(sdpb_inst_92_dout[29]),
  .I1(sdpb_inst_93_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1842 (
  .O(mux_o_1842),
  .I0(sdpb_inst_94_dout[29]),
  .I1(sdpb_inst_95_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1843 (
  .O(mux_o_1843),
  .I0(sdpb_inst_96_dout[29]),
  .I1(sdpb_inst_97_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1844 (
  .O(mux_o_1844),
  .I0(sdpb_inst_98_dout[29]),
  .I1(sdpb_inst_99_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1845 (
  .O(mux_o_1845),
  .I0(sdpb_inst_100_dout[29]),
  .I1(sdpb_inst_101_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1846 (
  .O(mux_o_1846),
  .I0(sdpb_inst_102_dout[29]),
  .I1(sdpb_inst_103_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1847 (
  .O(mux_o_1847),
  .I0(sdpb_inst_104_dout[29]),
  .I1(sdpb_inst_105_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1848 (
  .O(mux_o_1848),
  .I0(sdpb_inst_106_dout[29]),
  .I1(sdpb_inst_107_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1849 (
  .O(mux_o_1849),
  .I0(sdpb_inst_108_dout[29]),
  .I1(sdpb_inst_109_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1850 (
  .O(mux_o_1850),
  .I0(sdpb_inst_110_dout[29]),
  .I1(sdpb_inst_111_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1851 (
  .O(mux_o_1851),
  .I0(sdpb_inst_112_dout[29]),
  .I1(sdpb_inst_113_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1852 (
  .O(mux_o_1852),
  .I0(sdpb_inst_114_dout[29]),
  .I1(sdpb_inst_115_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1853 (
  .O(mux_o_1853),
  .I0(sdpb_inst_116_dout[29]),
  .I1(sdpb_inst_117_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1854 (
  .O(mux_o_1854),
  .I0(sdpb_inst_118_dout[29]),
  .I1(sdpb_inst_119_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1855 (
  .O(mux_o_1855),
  .I0(sdpb_inst_120_dout[29]),
  .I1(sdpb_inst_121_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1856 (
  .O(mux_o_1856),
  .I0(sdpb_inst_122_dout[29]),
  .I1(sdpb_inst_123_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1857 (
  .O(mux_o_1857),
  .I0(sdpb_inst_124_dout[29]),
  .I1(sdpb_inst_125_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1858 (
  .O(mux_o_1858),
  .I0(sdpb_inst_126_dout[29]),
  .I1(sdpb_inst_127_dout[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1859 (
  .O(mux_o_1859),
  .I0(mux_o_1827),
  .I1(mux_o_1828),
  .S0(dff_q_4)
);
MUX2 mux_inst_1860 (
  .O(mux_o_1860),
  .I0(mux_o_1829),
  .I1(mux_o_1830),
  .S0(dff_q_4)
);
MUX2 mux_inst_1861 (
  .O(mux_o_1861),
  .I0(mux_o_1831),
  .I1(mux_o_1832),
  .S0(dff_q_4)
);
MUX2 mux_inst_1862 (
  .O(mux_o_1862),
  .I0(mux_o_1833),
  .I1(mux_o_1834),
  .S0(dff_q_4)
);
MUX2 mux_inst_1863 (
  .O(mux_o_1863),
  .I0(mux_o_1835),
  .I1(mux_o_1836),
  .S0(dff_q_4)
);
MUX2 mux_inst_1864 (
  .O(mux_o_1864),
  .I0(mux_o_1837),
  .I1(mux_o_1838),
  .S0(dff_q_4)
);
MUX2 mux_inst_1865 (
  .O(mux_o_1865),
  .I0(mux_o_1839),
  .I1(mux_o_1840),
  .S0(dff_q_4)
);
MUX2 mux_inst_1866 (
  .O(mux_o_1866),
  .I0(mux_o_1841),
  .I1(mux_o_1842),
  .S0(dff_q_4)
);
MUX2 mux_inst_1867 (
  .O(mux_o_1867),
  .I0(mux_o_1843),
  .I1(mux_o_1844),
  .S0(dff_q_4)
);
MUX2 mux_inst_1868 (
  .O(mux_o_1868),
  .I0(mux_o_1845),
  .I1(mux_o_1846),
  .S0(dff_q_4)
);
MUX2 mux_inst_1869 (
  .O(mux_o_1869),
  .I0(mux_o_1847),
  .I1(mux_o_1848),
  .S0(dff_q_4)
);
MUX2 mux_inst_1870 (
  .O(mux_o_1870),
  .I0(mux_o_1849),
  .I1(mux_o_1850),
  .S0(dff_q_4)
);
MUX2 mux_inst_1871 (
  .O(mux_o_1871),
  .I0(mux_o_1851),
  .I1(mux_o_1852),
  .S0(dff_q_4)
);
MUX2 mux_inst_1872 (
  .O(mux_o_1872),
  .I0(mux_o_1853),
  .I1(mux_o_1854),
  .S0(dff_q_4)
);
MUX2 mux_inst_1873 (
  .O(mux_o_1873),
  .I0(mux_o_1855),
  .I1(mux_o_1856),
  .S0(dff_q_4)
);
MUX2 mux_inst_1874 (
  .O(mux_o_1874),
  .I0(mux_o_1857),
  .I1(mux_o_1858),
  .S0(dff_q_4)
);
MUX2 mux_inst_1875 (
  .O(mux_o_1875),
  .I0(mux_o_1859),
  .I1(mux_o_1860),
  .S0(dff_q_3)
);
MUX2 mux_inst_1876 (
  .O(mux_o_1876),
  .I0(mux_o_1861),
  .I1(mux_o_1862),
  .S0(dff_q_3)
);
MUX2 mux_inst_1877 (
  .O(mux_o_1877),
  .I0(mux_o_1863),
  .I1(mux_o_1864),
  .S0(dff_q_3)
);
MUX2 mux_inst_1878 (
  .O(mux_o_1878),
  .I0(mux_o_1865),
  .I1(mux_o_1866),
  .S0(dff_q_3)
);
MUX2 mux_inst_1879 (
  .O(mux_o_1879),
  .I0(mux_o_1867),
  .I1(mux_o_1868),
  .S0(dff_q_3)
);
MUX2 mux_inst_1880 (
  .O(mux_o_1880),
  .I0(mux_o_1869),
  .I1(mux_o_1870),
  .S0(dff_q_3)
);
MUX2 mux_inst_1881 (
  .O(mux_o_1881),
  .I0(mux_o_1871),
  .I1(mux_o_1872),
  .S0(dff_q_3)
);
MUX2 mux_inst_1882 (
  .O(mux_o_1882),
  .I0(mux_o_1873),
  .I1(mux_o_1874),
  .S0(dff_q_3)
);
MUX2 mux_inst_1883 (
  .O(mux_o_1883),
  .I0(mux_o_1875),
  .I1(mux_o_1876),
  .S0(dff_q_2)
);
MUX2 mux_inst_1884 (
  .O(mux_o_1884),
  .I0(mux_o_1877),
  .I1(mux_o_1878),
  .S0(dff_q_2)
);
MUX2 mux_inst_1885 (
  .O(mux_o_1885),
  .I0(mux_o_1879),
  .I1(mux_o_1880),
  .S0(dff_q_2)
);
MUX2 mux_inst_1886 (
  .O(mux_o_1886),
  .I0(mux_o_1881),
  .I1(mux_o_1882),
  .S0(dff_q_2)
);
MUX2 mux_inst_1887 (
  .O(mux_o_1887),
  .I0(mux_o_1883),
  .I1(mux_o_1884),
  .S0(dff_q_1)
);
MUX2 mux_inst_1888 (
  .O(mux_o_1888),
  .I0(mux_o_1885),
  .I1(mux_o_1886),
  .S0(dff_q_1)
);
MUX2 mux_inst_1889 (
  .O(dout[29]),
  .I0(mux_o_1887),
  .I1(mux_o_1888),
  .S0(dff_q_0)
);
MUX2 mux_inst_1890 (
  .O(mux_o_1890),
  .I0(sdpb_inst_64_dout[30]),
  .I1(sdpb_inst_65_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1891 (
  .O(mux_o_1891),
  .I0(sdpb_inst_66_dout[30]),
  .I1(sdpb_inst_67_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1892 (
  .O(mux_o_1892),
  .I0(sdpb_inst_68_dout[30]),
  .I1(sdpb_inst_69_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1893 (
  .O(mux_o_1893),
  .I0(sdpb_inst_70_dout[30]),
  .I1(sdpb_inst_71_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1894 (
  .O(mux_o_1894),
  .I0(sdpb_inst_72_dout[30]),
  .I1(sdpb_inst_73_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1895 (
  .O(mux_o_1895),
  .I0(sdpb_inst_74_dout[30]),
  .I1(sdpb_inst_75_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1896 (
  .O(mux_o_1896),
  .I0(sdpb_inst_76_dout[30]),
  .I1(sdpb_inst_77_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1897 (
  .O(mux_o_1897),
  .I0(sdpb_inst_78_dout[30]),
  .I1(sdpb_inst_79_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1898 (
  .O(mux_o_1898),
  .I0(sdpb_inst_80_dout[30]),
  .I1(sdpb_inst_81_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1899 (
  .O(mux_o_1899),
  .I0(sdpb_inst_82_dout[30]),
  .I1(sdpb_inst_83_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1900 (
  .O(mux_o_1900),
  .I0(sdpb_inst_84_dout[30]),
  .I1(sdpb_inst_85_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1901 (
  .O(mux_o_1901),
  .I0(sdpb_inst_86_dout[30]),
  .I1(sdpb_inst_87_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1902 (
  .O(mux_o_1902),
  .I0(sdpb_inst_88_dout[30]),
  .I1(sdpb_inst_89_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1903 (
  .O(mux_o_1903),
  .I0(sdpb_inst_90_dout[30]),
  .I1(sdpb_inst_91_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1904 (
  .O(mux_o_1904),
  .I0(sdpb_inst_92_dout[30]),
  .I1(sdpb_inst_93_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1905 (
  .O(mux_o_1905),
  .I0(sdpb_inst_94_dout[30]),
  .I1(sdpb_inst_95_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1906 (
  .O(mux_o_1906),
  .I0(sdpb_inst_96_dout[30]),
  .I1(sdpb_inst_97_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1907 (
  .O(mux_o_1907),
  .I0(sdpb_inst_98_dout[30]),
  .I1(sdpb_inst_99_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1908 (
  .O(mux_o_1908),
  .I0(sdpb_inst_100_dout[30]),
  .I1(sdpb_inst_101_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1909 (
  .O(mux_o_1909),
  .I0(sdpb_inst_102_dout[30]),
  .I1(sdpb_inst_103_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1910 (
  .O(mux_o_1910),
  .I0(sdpb_inst_104_dout[30]),
  .I1(sdpb_inst_105_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1911 (
  .O(mux_o_1911),
  .I0(sdpb_inst_106_dout[30]),
  .I1(sdpb_inst_107_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1912 (
  .O(mux_o_1912),
  .I0(sdpb_inst_108_dout[30]),
  .I1(sdpb_inst_109_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1913 (
  .O(mux_o_1913),
  .I0(sdpb_inst_110_dout[30]),
  .I1(sdpb_inst_111_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1914 (
  .O(mux_o_1914),
  .I0(sdpb_inst_112_dout[30]),
  .I1(sdpb_inst_113_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1915 (
  .O(mux_o_1915),
  .I0(sdpb_inst_114_dout[30]),
  .I1(sdpb_inst_115_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1916 (
  .O(mux_o_1916),
  .I0(sdpb_inst_116_dout[30]),
  .I1(sdpb_inst_117_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1917 (
  .O(mux_o_1917),
  .I0(sdpb_inst_118_dout[30]),
  .I1(sdpb_inst_119_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1918 (
  .O(mux_o_1918),
  .I0(sdpb_inst_120_dout[30]),
  .I1(sdpb_inst_121_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1919 (
  .O(mux_o_1919),
  .I0(sdpb_inst_122_dout[30]),
  .I1(sdpb_inst_123_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1920 (
  .O(mux_o_1920),
  .I0(sdpb_inst_124_dout[30]),
  .I1(sdpb_inst_125_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1921 (
  .O(mux_o_1921),
  .I0(sdpb_inst_126_dout[30]),
  .I1(sdpb_inst_127_dout[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1922 (
  .O(mux_o_1922),
  .I0(mux_o_1890),
  .I1(mux_o_1891),
  .S0(dff_q_4)
);
MUX2 mux_inst_1923 (
  .O(mux_o_1923),
  .I0(mux_o_1892),
  .I1(mux_o_1893),
  .S0(dff_q_4)
);
MUX2 mux_inst_1924 (
  .O(mux_o_1924),
  .I0(mux_o_1894),
  .I1(mux_o_1895),
  .S0(dff_q_4)
);
MUX2 mux_inst_1925 (
  .O(mux_o_1925),
  .I0(mux_o_1896),
  .I1(mux_o_1897),
  .S0(dff_q_4)
);
MUX2 mux_inst_1926 (
  .O(mux_o_1926),
  .I0(mux_o_1898),
  .I1(mux_o_1899),
  .S0(dff_q_4)
);
MUX2 mux_inst_1927 (
  .O(mux_o_1927),
  .I0(mux_o_1900),
  .I1(mux_o_1901),
  .S0(dff_q_4)
);
MUX2 mux_inst_1928 (
  .O(mux_o_1928),
  .I0(mux_o_1902),
  .I1(mux_o_1903),
  .S0(dff_q_4)
);
MUX2 mux_inst_1929 (
  .O(mux_o_1929),
  .I0(mux_o_1904),
  .I1(mux_o_1905),
  .S0(dff_q_4)
);
MUX2 mux_inst_1930 (
  .O(mux_o_1930),
  .I0(mux_o_1906),
  .I1(mux_o_1907),
  .S0(dff_q_4)
);
MUX2 mux_inst_1931 (
  .O(mux_o_1931),
  .I0(mux_o_1908),
  .I1(mux_o_1909),
  .S0(dff_q_4)
);
MUX2 mux_inst_1932 (
  .O(mux_o_1932),
  .I0(mux_o_1910),
  .I1(mux_o_1911),
  .S0(dff_q_4)
);
MUX2 mux_inst_1933 (
  .O(mux_o_1933),
  .I0(mux_o_1912),
  .I1(mux_o_1913),
  .S0(dff_q_4)
);
MUX2 mux_inst_1934 (
  .O(mux_o_1934),
  .I0(mux_o_1914),
  .I1(mux_o_1915),
  .S0(dff_q_4)
);
MUX2 mux_inst_1935 (
  .O(mux_o_1935),
  .I0(mux_o_1916),
  .I1(mux_o_1917),
  .S0(dff_q_4)
);
MUX2 mux_inst_1936 (
  .O(mux_o_1936),
  .I0(mux_o_1918),
  .I1(mux_o_1919),
  .S0(dff_q_4)
);
MUX2 mux_inst_1937 (
  .O(mux_o_1937),
  .I0(mux_o_1920),
  .I1(mux_o_1921),
  .S0(dff_q_4)
);
MUX2 mux_inst_1938 (
  .O(mux_o_1938),
  .I0(mux_o_1922),
  .I1(mux_o_1923),
  .S0(dff_q_3)
);
MUX2 mux_inst_1939 (
  .O(mux_o_1939),
  .I0(mux_o_1924),
  .I1(mux_o_1925),
  .S0(dff_q_3)
);
MUX2 mux_inst_1940 (
  .O(mux_o_1940),
  .I0(mux_o_1926),
  .I1(mux_o_1927),
  .S0(dff_q_3)
);
MUX2 mux_inst_1941 (
  .O(mux_o_1941),
  .I0(mux_o_1928),
  .I1(mux_o_1929),
  .S0(dff_q_3)
);
MUX2 mux_inst_1942 (
  .O(mux_o_1942),
  .I0(mux_o_1930),
  .I1(mux_o_1931),
  .S0(dff_q_3)
);
MUX2 mux_inst_1943 (
  .O(mux_o_1943),
  .I0(mux_o_1932),
  .I1(mux_o_1933),
  .S0(dff_q_3)
);
MUX2 mux_inst_1944 (
  .O(mux_o_1944),
  .I0(mux_o_1934),
  .I1(mux_o_1935),
  .S0(dff_q_3)
);
MUX2 mux_inst_1945 (
  .O(mux_o_1945),
  .I0(mux_o_1936),
  .I1(mux_o_1937),
  .S0(dff_q_3)
);
MUX2 mux_inst_1946 (
  .O(mux_o_1946),
  .I0(mux_o_1938),
  .I1(mux_o_1939),
  .S0(dff_q_2)
);
MUX2 mux_inst_1947 (
  .O(mux_o_1947),
  .I0(mux_o_1940),
  .I1(mux_o_1941),
  .S0(dff_q_2)
);
MUX2 mux_inst_1948 (
  .O(mux_o_1948),
  .I0(mux_o_1942),
  .I1(mux_o_1943),
  .S0(dff_q_2)
);
MUX2 mux_inst_1949 (
  .O(mux_o_1949),
  .I0(mux_o_1944),
  .I1(mux_o_1945),
  .S0(dff_q_2)
);
MUX2 mux_inst_1950 (
  .O(mux_o_1950),
  .I0(mux_o_1946),
  .I1(mux_o_1947),
  .S0(dff_q_1)
);
MUX2 mux_inst_1951 (
  .O(mux_o_1951),
  .I0(mux_o_1948),
  .I1(mux_o_1949),
  .S0(dff_q_1)
);
MUX2 mux_inst_1952 (
  .O(dout[30]),
  .I0(mux_o_1950),
  .I1(mux_o_1951),
  .S0(dff_q_0)
);
MUX2 mux_inst_1953 (
  .O(mux_o_1953),
  .I0(sdpb_inst_64_dout[31]),
  .I1(sdpb_inst_65_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1954 (
  .O(mux_o_1954),
  .I0(sdpb_inst_66_dout[31]),
  .I1(sdpb_inst_67_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1955 (
  .O(mux_o_1955),
  .I0(sdpb_inst_68_dout[31]),
  .I1(sdpb_inst_69_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1956 (
  .O(mux_o_1956),
  .I0(sdpb_inst_70_dout[31]),
  .I1(sdpb_inst_71_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1957 (
  .O(mux_o_1957),
  .I0(sdpb_inst_72_dout[31]),
  .I1(sdpb_inst_73_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1958 (
  .O(mux_o_1958),
  .I0(sdpb_inst_74_dout[31]),
  .I1(sdpb_inst_75_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1959 (
  .O(mux_o_1959),
  .I0(sdpb_inst_76_dout[31]),
  .I1(sdpb_inst_77_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1960 (
  .O(mux_o_1960),
  .I0(sdpb_inst_78_dout[31]),
  .I1(sdpb_inst_79_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1961 (
  .O(mux_o_1961),
  .I0(sdpb_inst_80_dout[31]),
  .I1(sdpb_inst_81_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1962 (
  .O(mux_o_1962),
  .I0(sdpb_inst_82_dout[31]),
  .I1(sdpb_inst_83_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1963 (
  .O(mux_o_1963),
  .I0(sdpb_inst_84_dout[31]),
  .I1(sdpb_inst_85_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1964 (
  .O(mux_o_1964),
  .I0(sdpb_inst_86_dout[31]),
  .I1(sdpb_inst_87_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1965 (
  .O(mux_o_1965),
  .I0(sdpb_inst_88_dout[31]),
  .I1(sdpb_inst_89_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1966 (
  .O(mux_o_1966),
  .I0(sdpb_inst_90_dout[31]),
  .I1(sdpb_inst_91_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1967 (
  .O(mux_o_1967),
  .I0(sdpb_inst_92_dout[31]),
  .I1(sdpb_inst_93_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1968 (
  .O(mux_o_1968),
  .I0(sdpb_inst_94_dout[31]),
  .I1(sdpb_inst_95_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1969 (
  .O(mux_o_1969),
  .I0(sdpb_inst_96_dout[31]),
  .I1(sdpb_inst_97_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1970 (
  .O(mux_o_1970),
  .I0(sdpb_inst_98_dout[31]),
  .I1(sdpb_inst_99_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1971 (
  .O(mux_o_1971),
  .I0(sdpb_inst_100_dout[31]),
  .I1(sdpb_inst_101_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1972 (
  .O(mux_o_1972),
  .I0(sdpb_inst_102_dout[31]),
  .I1(sdpb_inst_103_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1973 (
  .O(mux_o_1973),
  .I0(sdpb_inst_104_dout[31]),
  .I1(sdpb_inst_105_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1974 (
  .O(mux_o_1974),
  .I0(sdpb_inst_106_dout[31]),
  .I1(sdpb_inst_107_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1975 (
  .O(mux_o_1975),
  .I0(sdpb_inst_108_dout[31]),
  .I1(sdpb_inst_109_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1976 (
  .O(mux_o_1976),
  .I0(sdpb_inst_110_dout[31]),
  .I1(sdpb_inst_111_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1977 (
  .O(mux_o_1977),
  .I0(sdpb_inst_112_dout[31]),
  .I1(sdpb_inst_113_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1978 (
  .O(mux_o_1978),
  .I0(sdpb_inst_114_dout[31]),
  .I1(sdpb_inst_115_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1979 (
  .O(mux_o_1979),
  .I0(sdpb_inst_116_dout[31]),
  .I1(sdpb_inst_117_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1980 (
  .O(mux_o_1980),
  .I0(sdpb_inst_118_dout[31]),
  .I1(sdpb_inst_119_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1981 (
  .O(mux_o_1981),
  .I0(sdpb_inst_120_dout[31]),
  .I1(sdpb_inst_121_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1982 (
  .O(mux_o_1982),
  .I0(sdpb_inst_122_dout[31]),
  .I1(sdpb_inst_123_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1983 (
  .O(mux_o_1983),
  .I0(sdpb_inst_124_dout[31]),
  .I1(sdpb_inst_125_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1984 (
  .O(mux_o_1984),
  .I0(sdpb_inst_126_dout[31]),
  .I1(sdpb_inst_127_dout[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1985 (
  .O(mux_o_1985),
  .I0(mux_o_1953),
  .I1(mux_o_1954),
  .S0(dff_q_4)
);
MUX2 mux_inst_1986 (
  .O(mux_o_1986),
  .I0(mux_o_1955),
  .I1(mux_o_1956),
  .S0(dff_q_4)
);
MUX2 mux_inst_1987 (
  .O(mux_o_1987),
  .I0(mux_o_1957),
  .I1(mux_o_1958),
  .S0(dff_q_4)
);
MUX2 mux_inst_1988 (
  .O(mux_o_1988),
  .I0(mux_o_1959),
  .I1(mux_o_1960),
  .S0(dff_q_4)
);
MUX2 mux_inst_1989 (
  .O(mux_o_1989),
  .I0(mux_o_1961),
  .I1(mux_o_1962),
  .S0(dff_q_4)
);
MUX2 mux_inst_1990 (
  .O(mux_o_1990),
  .I0(mux_o_1963),
  .I1(mux_o_1964),
  .S0(dff_q_4)
);
MUX2 mux_inst_1991 (
  .O(mux_o_1991),
  .I0(mux_o_1965),
  .I1(mux_o_1966),
  .S0(dff_q_4)
);
MUX2 mux_inst_1992 (
  .O(mux_o_1992),
  .I0(mux_o_1967),
  .I1(mux_o_1968),
  .S0(dff_q_4)
);
MUX2 mux_inst_1993 (
  .O(mux_o_1993),
  .I0(mux_o_1969),
  .I1(mux_o_1970),
  .S0(dff_q_4)
);
MUX2 mux_inst_1994 (
  .O(mux_o_1994),
  .I0(mux_o_1971),
  .I1(mux_o_1972),
  .S0(dff_q_4)
);
MUX2 mux_inst_1995 (
  .O(mux_o_1995),
  .I0(mux_o_1973),
  .I1(mux_o_1974),
  .S0(dff_q_4)
);
MUX2 mux_inst_1996 (
  .O(mux_o_1996),
  .I0(mux_o_1975),
  .I1(mux_o_1976),
  .S0(dff_q_4)
);
MUX2 mux_inst_1997 (
  .O(mux_o_1997),
  .I0(mux_o_1977),
  .I1(mux_o_1978),
  .S0(dff_q_4)
);
MUX2 mux_inst_1998 (
  .O(mux_o_1998),
  .I0(mux_o_1979),
  .I1(mux_o_1980),
  .S0(dff_q_4)
);
MUX2 mux_inst_1999 (
  .O(mux_o_1999),
  .I0(mux_o_1981),
  .I1(mux_o_1982),
  .S0(dff_q_4)
);
MUX2 mux_inst_2000 (
  .O(mux_o_2000),
  .I0(mux_o_1983),
  .I1(mux_o_1984),
  .S0(dff_q_4)
);
MUX2 mux_inst_2001 (
  .O(mux_o_2001),
  .I0(mux_o_1985),
  .I1(mux_o_1986),
  .S0(dff_q_3)
);
MUX2 mux_inst_2002 (
  .O(mux_o_2002),
  .I0(mux_o_1987),
  .I1(mux_o_1988),
  .S0(dff_q_3)
);
MUX2 mux_inst_2003 (
  .O(mux_o_2003),
  .I0(mux_o_1989),
  .I1(mux_o_1990),
  .S0(dff_q_3)
);
MUX2 mux_inst_2004 (
  .O(mux_o_2004),
  .I0(mux_o_1991),
  .I1(mux_o_1992),
  .S0(dff_q_3)
);
MUX2 mux_inst_2005 (
  .O(mux_o_2005),
  .I0(mux_o_1993),
  .I1(mux_o_1994),
  .S0(dff_q_3)
);
MUX2 mux_inst_2006 (
  .O(mux_o_2006),
  .I0(mux_o_1995),
  .I1(mux_o_1996),
  .S0(dff_q_3)
);
MUX2 mux_inst_2007 (
  .O(mux_o_2007),
  .I0(mux_o_1997),
  .I1(mux_o_1998),
  .S0(dff_q_3)
);
MUX2 mux_inst_2008 (
  .O(mux_o_2008),
  .I0(mux_o_1999),
  .I1(mux_o_2000),
  .S0(dff_q_3)
);
MUX2 mux_inst_2009 (
  .O(mux_o_2009),
  .I0(mux_o_2001),
  .I1(mux_o_2002),
  .S0(dff_q_2)
);
MUX2 mux_inst_2010 (
  .O(mux_o_2010),
  .I0(mux_o_2003),
  .I1(mux_o_2004),
  .S0(dff_q_2)
);
MUX2 mux_inst_2011 (
  .O(mux_o_2011),
  .I0(mux_o_2005),
  .I1(mux_o_2006),
  .S0(dff_q_2)
);
MUX2 mux_inst_2012 (
  .O(mux_o_2012),
  .I0(mux_o_2007),
  .I1(mux_o_2008),
  .S0(dff_q_2)
);
MUX2 mux_inst_2013 (
  .O(mux_o_2013),
  .I0(mux_o_2009),
  .I1(mux_o_2010),
  .S0(dff_q_1)
);
MUX2 mux_inst_2014 (
  .O(mux_o_2014),
  .I0(mux_o_2011),
  .I1(mux_o_2012),
  .S0(dff_q_1)
);
MUX2 mux_inst_2015 (
  .O(dout[31]),
  .I0(mux_o_2013),
  .I1(mux_o_2014),
  .S0(dff_q_0)
);
endmodule //SRAM_SDPB
