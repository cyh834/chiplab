module gw_gao(
    \asic/cpu/cpu/if_stage/fs_pc[31] ,
    \asic/cpu/cpu/if_stage/fs_pc[30] ,
    \asic/cpu/cpu/if_stage/fs_pc[29] ,
    \asic/cpu/cpu/if_stage/fs_pc[28] ,
    \asic/cpu/cpu/if_stage/fs_pc[27] ,
    \asic/cpu/cpu/if_stage/fs_pc[26] ,
    \asic/cpu/cpu/if_stage/fs_pc[25] ,
    \asic/cpu/cpu/if_stage/fs_pc[24] ,
    \asic/cpu/cpu/if_stage/fs_pc[23] ,
    \asic/cpu/cpu/if_stage/fs_pc[22] ,
    \asic/cpu/cpu/if_stage/fs_pc[21] ,
    \asic/cpu/cpu/if_stage/fs_pc[20] ,
    \asic/cpu/cpu/if_stage/fs_pc[19] ,
    \asic/cpu/cpu/if_stage/fs_pc[18] ,
    \asic/cpu/cpu/if_stage/fs_pc[17] ,
    \asic/cpu/cpu/if_stage/fs_pc[16] ,
    \asic/cpu/cpu/if_stage/fs_pc[15] ,
    \asic/cpu/cpu/if_stage/fs_pc[14] ,
    \asic/cpu/cpu/if_stage/fs_pc[13] ,
    \asic/cpu/cpu/if_stage/fs_pc[12] ,
    \asic/cpu/cpu/if_stage/fs_pc[11] ,
    \asic/cpu/cpu/if_stage/fs_pc[10] ,
    \asic/cpu/cpu/if_stage/fs_pc[9] ,
    \asic/cpu/cpu/if_stage/fs_pc[8] ,
    \asic/cpu/cpu/if_stage/fs_pc[7] ,
    \asic/cpu/cpu/if_stage/fs_pc[6] ,
    \asic/cpu/cpu/if_stage/fs_pc[5] ,
    \asic/cpu/cpu/if_stage/fs_pc[4] ,
    \asic/cpu/cpu/if_stage/fs_pc[3] ,
    \asic/cpu/cpu/if_stage/fs_pc[2] ,
    \asic/cpu/cpu/if_stage/fs_pc[1] ,
    \asic/cpu/cpu/if_stage/fs_pc[0] ,
    \asic/cpu/cpu/if_stage/fs_inst[31] ,
    \asic/cpu/cpu/if_stage/fs_inst[30] ,
    \asic/cpu/cpu/if_stage/fs_inst[29] ,
    \asic/cpu/cpu/if_stage/fs_inst[28] ,
    \asic/cpu/cpu/if_stage/fs_inst[27] ,
    \asic/cpu/cpu/if_stage/fs_inst[26] ,
    \asic/cpu/cpu/if_stage/fs_inst[25] ,
    \asic/cpu/cpu/if_stage/fs_inst[24] ,
    \asic/cpu/cpu/if_stage/fs_inst[23] ,
    \asic/cpu/cpu/if_stage/fs_inst[22] ,
    \asic/cpu/cpu/if_stage/fs_inst[21] ,
    \asic/cpu/cpu/if_stage/fs_inst[20] ,
    \asic/cpu/cpu/if_stage/fs_inst[19] ,
    \asic/cpu/cpu/if_stage/fs_inst[18] ,
    \asic/cpu/cpu/if_stage/fs_inst[17] ,
    \asic/cpu/cpu/if_stage/fs_inst[16] ,
    \asic/cpu/cpu/if_stage/fs_inst[15] ,
    \asic/cpu/cpu/if_stage/fs_inst[14] ,
    \asic/cpu/cpu/if_stage/fs_inst[13] ,
    \asic/cpu/cpu/if_stage/fs_inst[12] ,
    \asic/cpu/cpu/if_stage/fs_inst[11] ,
    \asic/cpu/cpu/if_stage/fs_inst[10] ,
    \asic/cpu/cpu/if_stage/fs_inst[9] ,
    \asic/cpu/cpu/if_stage/fs_inst[8] ,
    \asic/cpu/cpu/if_stage/fs_inst[7] ,
    \asic/cpu/cpu/if_stage/fs_inst[6] ,
    \asic/cpu/cpu/if_stage/fs_inst[5] ,
    \asic/cpu/cpu/if_stage/fs_inst[4] ,
    \asic/cpu/cpu/if_stage/fs_inst[3] ,
    \asic/cpu/cpu/if_stage/fs_inst[2] ,
    \asic/cpu/cpu/if_stage/fs_inst[1] ,
    \asic/cpu/cpu/if_stage/fs_inst[0] ,
    \asic/lsdram/msdram/io_in_awid[3] ,
    \asic/lsdram/msdram/io_in_awid[2] ,
    \asic/lsdram/msdram/io_in_awid[1] ,
    \asic/lsdram/msdram/io_in_awid[0] ,
    \asic/lsdram/msdram/io_in_awaddr[31] ,
    \asic/lsdram/msdram/io_in_awaddr[30] ,
    \asic/lsdram/msdram/io_in_awaddr[29] ,
    \asic/lsdram/msdram/io_in_awaddr[28] ,
    \asic/lsdram/msdram/io_in_awaddr[27] ,
    \asic/lsdram/msdram/io_in_awaddr[26] ,
    \asic/lsdram/msdram/io_in_awaddr[25] ,
    \asic/lsdram/msdram/io_in_awaddr[24] ,
    \asic/lsdram/msdram/io_in_awaddr[23] ,
    \asic/lsdram/msdram/io_in_awaddr[22] ,
    \asic/lsdram/msdram/io_in_awaddr[21] ,
    \asic/lsdram/msdram/io_in_awaddr[20] ,
    \asic/lsdram/msdram/io_in_awaddr[19] ,
    \asic/lsdram/msdram/io_in_awaddr[18] ,
    \asic/lsdram/msdram/io_in_awaddr[17] ,
    \asic/lsdram/msdram/io_in_awaddr[16] ,
    \asic/lsdram/msdram/io_in_awaddr[15] ,
    \asic/lsdram/msdram/io_in_awaddr[14] ,
    \asic/lsdram/msdram/io_in_awaddr[13] ,
    \asic/lsdram/msdram/io_in_awaddr[12] ,
    \asic/lsdram/msdram/io_in_awaddr[11] ,
    \asic/lsdram/msdram/io_in_awaddr[10] ,
    \asic/lsdram/msdram/io_in_awaddr[9] ,
    \asic/lsdram/msdram/io_in_awaddr[8] ,
    \asic/lsdram/msdram/io_in_awaddr[7] ,
    \asic/lsdram/msdram/io_in_awaddr[6] ,
    \asic/lsdram/msdram/io_in_awaddr[5] ,
    \asic/lsdram/msdram/io_in_awaddr[4] ,
    \asic/lsdram/msdram/io_in_awaddr[3] ,
    \asic/lsdram/msdram/io_in_awaddr[2] ,
    \asic/lsdram/msdram/io_in_awaddr[1] ,
    \asic/lsdram/msdram/io_in_awaddr[0] ,
    \asic/lsdram/msdram/io_in_awlen[7] ,
    \asic/lsdram/msdram/io_in_awlen[6] ,
    \asic/lsdram/msdram/io_in_awlen[5] ,
    \asic/lsdram/msdram/io_in_awlen[4] ,
    \asic/lsdram/msdram/io_in_awlen[3] ,
    \asic/lsdram/msdram/io_in_awlen[2] ,
    \asic/lsdram/msdram/io_in_awlen[1] ,
    \asic/lsdram/msdram/io_in_awlen[0] ,
    \asic/lsdram/msdram/io_in_awsize[2] ,
    \asic/lsdram/msdram/io_in_awsize[1] ,
    \asic/lsdram/msdram/io_in_awsize[0] ,
    \asic/lsdram/msdram/io_in_wdata[31] ,
    \asic/lsdram/msdram/io_in_wdata[30] ,
    \asic/lsdram/msdram/io_in_wdata[29] ,
    \asic/lsdram/msdram/io_in_wdata[28] ,
    \asic/lsdram/msdram/io_in_wdata[27] ,
    \asic/lsdram/msdram/io_in_wdata[26] ,
    \asic/lsdram/msdram/io_in_wdata[25] ,
    \asic/lsdram/msdram/io_in_wdata[24] ,
    \asic/lsdram/msdram/io_in_wdata[23] ,
    \asic/lsdram/msdram/io_in_wdata[22] ,
    \asic/lsdram/msdram/io_in_wdata[21] ,
    \asic/lsdram/msdram/io_in_wdata[20] ,
    \asic/lsdram/msdram/io_in_wdata[19] ,
    \asic/lsdram/msdram/io_in_wdata[18] ,
    \asic/lsdram/msdram/io_in_wdata[17] ,
    \asic/lsdram/msdram/io_in_wdata[16] ,
    \asic/lsdram/msdram/io_in_wdata[15] ,
    \asic/lsdram/msdram/io_in_wdata[14] ,
    \asic/lsdram/msdram/io_in_wdata[13] ,
    \asic/lsdram/msdram/io_in_wdata[12] ,
    \asic/lsdram/msdram/io_in_wdata[11] ,
    \asic/lsdram/msdram/io_in_wdata[10] ,
    \asic/lsdram/msdram/io_in_wdata[9] ,
    \asic/lsdram/msdram/io_in_wdata[8] ,
    \asic/lsdram/msdram/io_in_wdata[7] ,
    \asic/lsdram/msdram/io_in_wdata[6] ,
    \asic/lsdram/msdram/io_in_wdata[5] ,
    \asic/lsdram/msdram/io_in_wdata[4] ,
    \asic/lsdram/msdram/io_in_wdata[3] ,
    \asic/lsdram/msdram/io_in_wdata[2] ,
    \asic/lsdram/msdram/io_in_wdata[1] ,
    \asic/lsdram/msdram/io_in_wdata[0] ,
    \asic/lsdram/msdram/io_in_wstrb[3] ,
    \asic/lsdram/msdram/io_in_wstrb[2] ,
    \asic/lsdram/msdram/io_in_wstrb[1] ,
    \asic/lsdram/msdram/io_in_wstrb[0] ,
    \asic/lsdram/msdram/io_in_bid[3] ,
    \asic/lsdram/msdram/io_in_bid[2] ,
    \asic/lsdram/msdram/io_in_bid[1] ,
    \asic/lsdram/msdram/io_in_bid[0] ,
    \asic/lsdram/msdram/io_in_arid[3] ,
    \asic/lsdram/msdram/io_in_arid[2] ,
    \asic/lsdram/msdram/io_in_arid[1] ,
    \asic/lsdram/msdram/io_in_arid[0] ,
    \asic/lsdram/msdram/io_in_araddr[31] ,
    \asic/lsdram/msdram/io_in_araddr[30] ,
    \asic/lsdram/msdram/io_in_araddr[29] ,
    \asic/lsdram/msdram/io_in_araddr[28] ,
    \asic/lsdram/msdram/io_in_araddr[27] ,
    \asic/lsdram/msdram/io_in_araddr[26] ,
    \asic/lsdram/msdram/io_in_araddr[25] ,
    \asic/lsdram/msdram/io_in_araddr[24] ,
    \asic/lsdram/msdram/io_in_araddr[23] ,
    \asic/lsdram/msdram/io_in_araddr[22] ,
    \asic/lsdram/msdram/io_in_araddr[21] ,
    \asic/lsdram/msdram/io_in_araddr[20] ,
    \asic/lsdram/msdram/io_in_araddr[19] ,
    \asic/lsdram/msdram/io_in_araddr[18] ,
    \asic/lsdram/msdram/io_in_araddr[17] ,
    \asic/lsdram/msdram/io_in_araddr[16] ,
    \asic/lsdram/msdram/io_in_araddr[15] ,
    \asic/lsdram/msdram/io_in_araddr[14] ,
    \asic/lsdram/msdram/io_in_araddr[13] ,
    \asic/lsdram/msdram/io_in_araddr[12] ,
    \asic/lsdram/msdram/io_in_araddr[11] ,
    \asic/lsdram/msdram/io_in_araddr[10] ,
    \asic/lsdram/msdram/io_in_araddr[9] ,
    \asic/lsdram/msdram/io_in_araddr[8] ,
    \asic/lsdram/msdram/io_in_araddr[7] ,
    \asic/lsdram/msdram/io_in_araddr[6] ,
    \asic/lsdram/msdram/io_in_araddr[5] ,
    \asic/lsdram/msdram/io_in_araddr[4] ,
    \asic/lsdram/msdram/io_in_araddr[3] ,
    \asic/lsdram/msdram/io_in_araddr[2] ,
    \asic/lsdram/msdram/io_in_araddr[1] ,
    \asic/lsdram/msdram/io_in_araddr[0] ,
    \asic/lsdram/msdram/io_in_arlen[7] ,
    \asic/lsdram/msdram/io_in_arlen[6] ,
    \asic/lsdram/msdram/io_in_arlen[5] ,
    \asic/lsdram/msdram/io_in_arlen[4] ,
    \asic/lsdram/msdram/io_in_arlen[3] ,
    \asic/lsdram/msdram/io_in_arlen[2] ,
    \asic/lsdram/msdram/io_in_arlen[1] ,
    \asic/lsdram/msdram/io_in_arlen[0] ,
    \asic/lsdram/msdram/io_in_arsize[2] ,
    \asic/lsdram/msdram/io_in_arsize[1] ,
    \asic/lsdram/msdram/io_in_arsize[0] ,
    \asic/lsdram/msdram/io_in_rid[3] ,
    \asic/lsdram/msdram/io_in_rid[2] ,
    \asic/lsdram/msdram/io_in_rid[1] ,
    \asic/lsdram/msdram/io_in_rid[0] ,
    \asic/lsdram/msdram/io_in_rdata[31] ,
    \asic/lsdram/msdram/io_in_rdata[30] ,
    \asic/lsdram/msdram/io_in_rdata[29] ,
    \asic/lsdram/msdram/io_in_rdata[28] ,
    \asic/lsdram/msdram/io_in_rdata[27] ,
    \asic/lsdram/msdram/io_in_rdata[26] ,
    \asic/lsdram/msdram/io_in_rdata[25] ,
    \asic/lsdram/msdram/io_in_rdata[24] ,
    \asic/lsdram/msdram/io_in_rdata[23] ,
    \asic/lsdram/msdram/io_in_rdata[22] ,
    \asic/lsdram/msdram/io_in_rdata[21] ,
    \asic/lsdram/msdram/io_in_rdata[20] ,
    \asic/lsdram/msdram/io_in_rdata[19] ,
    \asic/lsdram/msdram/io_in_rdata[18] ,
    \asic/lsdram/msdram/io_in_rdata[17] ,
    \asic/lsdram/msdram/io_in_rdata[16] ,
    \asic/lsdram/msdram/io_in_rdata[15] ,
    \asic/lsdram/msdram/io_in_rdata[14] ,
    \asic/lsdram/msdram/io_in_rdata[13] ,
    \asic/lsdram/msdram/io_in_rdata[12] ,
    \asic/lsdram/msdram/io_in_rdata[11] ,
    \asic/lsdram/msdram/io_in_rdata[10] ,
    \asic/lsdram/msdram/io_in_rdata[9] ,
    \asic/lsdram/msdram/io_in_rdata[8] ,
    \asic/lsdram/msdram/io_in_rdata[7] ,
    \asic/lsdram/msdram/io_in_rdata[6] ,
    \asic/lsdram/msdram/io_in_rdata[5] ,
    \asic/lsdram/msdram/io_in_rdata[4] ,
    \asic/lsdram/msdram/io_in_rdata[3] ,
    \asic/lsdram/msdram/io_in_rdata[2] ,
    \asic/lsdram/msdram/io_in_rdata[1] ,
    \asic/lsdram/msdram/io_in_rdata[0] ,
    \asic/lsdram/msdram/io_dmi_cmd[2] ,
    \asic/lsdram/msdram/io_dmi_cmd[1] ,
    \asic/lsdram/msdram/io_dmi_cmd[0] ,
    \asic/lsdram/msdram/io_dmi_addr[28] ,
    \asic/lsdram/msdram/io_dmi_addr[27] ,
    \asic/lsdram/msdram/io_dmi_addr[26] ,
    \asic/lsdram/msdram/io_dmi_addr[25] ,
    \asic/lsdram/msdram/io_dmi_addr[24] ,
    \asic/lsdram/msdram/io_dmi_addr[23] ,
    \asic/lsdram/msdram/io_dmi_addr[22] ,
    \asic/lsdram/msdram/io_dmi_addr[21] ,
    \asic/lsdram/msdram/io_dmi_addr[20] ,
    \asic/lsdram/msdram/io_dmi_addr[19] ,
    \asic/lsdram/msdram/io_dmi_addr[18] ,
    \asic/lsdram/msdram/io_dmi_addr[17] ,
    \asic/lsdram/msdram/io_dmi_addr[16] ,
    \asic/lsdram/msdram/io_dmi_addr[15] ,
    \asic/lsdram/msdram/io_dmi_addr[14] ,
    \asic/lsdram/msdram/io_dmi_addr[13] ,
    \asic/lsdram/msdram/io_dmi_addr[12] ,
    \asic/lsdram/msdram/io_dmi_addr[11] ,
    \asic/lsdram/msdram/io_dmi_addr[10] ,
    \asic/lsdram/msdram/io_dmi_addr[9] ,
    \asic/lsdram/msdram/io_dmi_addr[8] ,
    \asic/lsdram/msdram/io_dmi_addr[7] ,
    \asic/lsdram/msdram/io_dmi_addr[6] ,
    \asic/lsdram/msdram/io_dmi_addr[5] ,
    \asic/lsdram/msdram/io_dmi_addr[4] ,
    \asic/lsdram/msdram/io_dmi_addr[3] ,
    \asic/lsdram/msdram/io_dmi_addr[2] ,
    \asic/lsdram/msdram/io_dmi_addr[1] ,
    \asic/lsdram/msdram/io_dmi_addr[0] ,
    \asic/lsdram/msdram/io_dmi_wr_data[255] ,
    \asic/lsdram/msdram/io_dmi_wr_data[254] ,
    \asic/lsdram/msdram/io_dmi_wr_data[253] ,
    \asic/lsdram/msdram/io_dmi_wr_data[252] ,
    \asic/lsdram/msdram/io_dmi_wr_data[251] ,
    \asic/lsdram/msdram/io_dmi_wr_data[250] ,
    \asic/lsdram/msdram/io_dmi_wr_data[249] ,
    \asic/lsdram/msdram/io_dmi_wr_data[248] ,
    \asic/lsdram/msdram/io_dmi_wr_data[247] ,
    \asic/lsdram/msdram/io_dmi_wr_data[246] ,
    \asic/lsdram/msdram/io_dmi_wr_data[245] ,
    \asic/lsdram/msdram/io_dmi_wr_data[244] ,
    \asic/lsdram/msdram/io_dmi_wr_data[243] ,
    \asic/lsdram/msdram/io_dmi_wr_data[242] ,
    \asic/lsdram/msdram/io_dmi_wr_data[241] ,
    \asic/lsdram/msdram/io_dmi_wr_data[240] ,
    \asic/lsdram/msdram/io_dmi_wr_data[239] ,
    \asic/lsdram/msdram/io_dmi_wr_data[238] ,
    \asic/lsdram/msdram/io_dmi_wr_data[237] ,
    \asic/lsdram/msdram/io_dmi_wr_data[236] ,
    \asic/lsdram/msdram/io_dmi_wr_data[235] ,
    \asic/lsdram/msdram/io_dmi_wr_data[234] ,
    \asic/lsdram/msdram/io_dmi_wr_data[233] ,
    \asic/lsdram/msdram/io_dmi_wr_data[232] ,
    \asic/lsdram/msdram/io_dmi_wr_data[231] ,
    \asic/lsdram/msdram/io_dmi_wr_data[230] ,
    \asic/lsdram/msdram/io_dmi_wr_data[229] ,
    \asic/lsdram/msdram/io_dmi_wr_data[228] ,
    \asic/lsdram/msdram/io_dmi_wr_data[227] ,
    \asic/lsdram/msdram/io_dmi_wr_data[226] ,
    \asic/lsdram/msdram/io_dmi_wr_data[225] ,
    \asic/lsdram/msdram/io_dmi_wr_data[224] ,
    \asic/lsdram/msdram/io_dmi_wr_data[223] ,
    \asic/lsdram/msdram/io_dmi_wr_data[222] ,
    \asic/lsdram/msdram/io_dmi_wr_data[221] ,
    \asic/lsdram/msdram/io_dmi_wr_data[220] ,
    \asic/lsdram/msdram/io_dmi_wr_data[219] ,
    \asic/lsdram/msdram/io_dmi_wr_data[218] ,
    \asic/lsdram/msdram/io_dmi_wr_data[217] ,
    \asic/lsdram/msdram/io_dmi_wr_data[216] ,
    \asic/lsdram/msdram/io_dmi_wr_data[215] ,
    \asic/lsdram/msdram/io_dmi_wr_data[214] ,
    \asic/lsdram/msdram/io_dmi_wr_data[213] ,
    \asic/lsdram/msdram/io_dmi_wr_data[212] ,
    \asic/lsdram/msdram/io_dmi_wr_data[211] ,
    \asic/lsdram/msdram/io_dmi_wr_data[210] ,
    \asic/lsdram/msdram/io_dmi_wr_data[209] ,
    \asic/lsdram/msdram/io_dmi_wr_data[208] ,
    \asic/lsdram/msdram/io_dmi_wr_data[207] ,
    \asic/lsdram/msdram/io_dmi_wr_data[206] ,
    \asic/lsdram/msdram/io_dmi_wr_data[205] ,
    \asic/lsdram/msdram/io_dmi_wr_data[204] ,
    \asic/lsdram/msdram/io_dmi_wr_data[203] ,
    \asic/lsdram/msdram/io_dmi_wr_data[202] ,
    \asic/lsdram/msdram/io_dmi_wr_data[201] ,
    \asic/lsdram/msdram/io_dmi_wr_data[200] ,
    \asic/lsdram/msdram/io_dmi_wr_data[199] ,
    \asic/lsdram/msdram/io_dmi_wr_data[198] ,
    \asic/lsdram/msdram/io_dmi_wr_data[197] ,
    \asic/lsdram/msdram/io_dmi_wr_data[196] ,
    \asic/lsdram/msdram/io_dmi_wr_data[195] ,
    \asic/lsdram/msdram/io_dmi_wr_data[194] ,
    \asic/lsdram/msdram/io_dmi_wr_data[193] ,
    \asic/lsdram/msdram/io_dmi_wr_data[192] ,
    \asic/lsdram/msdram/io_dmi_wr_data[191] ,
    \asic/lsdram/msdram/io_dmi_wr_data[190] ,
    \asic/lsdram/msdram/io_dmi_wr_data[189] ,
    \asic/lsdram/msdram/io_dmi_wr_data[188] ,
    \asic/lsdram/msdram/io_dmi_wr_data[187] ,
    \asic/lsdram/msdram/io_dmi_wr_data[186] ,
    \asic/lsdram/msdram/io_dmi_wr_data[185] ,
    \asic/lsdram/msdram/io_dmi_wr_data[184] ,
    \asic/lsdram/msdram/io_dmi_wr_data[183] ,
    \asic/lsdram/msdram/io_dmi_wr_data[182] ,
    \asic/lsdram/msdram/io_dmi_wr_data[181] ,
    \asic/lsdram/msdram/io_dmi_wr_data[180] ,
    \asic/lsdram/msdram/io_dmi_wr_data[179] ,
    \asic/lsdram/msdram/io_dmi_wr_data[178] ,
    \asic/lsdram/msdram/io_dmi_wr_data[177] ,
    \asic/lsdram/msdram/io_dmi_wr_data[176] ,
    \asic/lsdram/msdram/io_dmi_wr_data[175] ,
    \asic/lsdram/msdram/io_dmi_wr_data[174] ,
    \asic/lsdram/msdram/io_dmi_wr_data[173] ,
    \asic/lsdram/msdram/io_dmi_wr_data[172] ,
    \asic/lsdram/msdram/io_dmi_wr_data[171] ,
    \asic/lsdram/msdram/io_dmi_wr_data[170] ,
    \asic/lsdram/msdram/io_dmi_wr_data[169] ,
    \asic/lsdram/msdram/io_dmi_wr_data[168] ,
    \asic/lsdram/msdram/io_dmi_wr_data[167] ,
    \asic/lsdram/msdram/io_dmi_wr_data[166] ,
    \asic/lsdram/msdram/io_dmi_wr_data[165] ,
    \asic/lsdram/msdram/io_dmi_wr_data[164] ,
    \asic/lsdram/msdram/io_dmi_wr_data[163] ,
    \asic/lsdram/msdram/io_dmi_wr_data[162] ,
    \asic/lsdram/msdram/io_dmi_wr_data[161] ,
    \asic/lsdram/msdram/io_dmi_wr_data[160] ,
    \asic/lsdram/msdram/io_dmi_wr_data[159] ,
    \asic/lsdram/msdram/io_dmi_wr_data[158] ,
    \asic/lsdram/msdram/io_dmi_wr_data[157] ,
    \asic/lsdram/msdram/io_dmi_wr_data[156] ,
    \asic/lsdram/msdram/io_dmi_wr_data[155] ,
    \asic/lsdram/msdram/io_dmi_wr_data[154] ,
    \asic/lsdram/msdram/io_dmi_wr_data[153] ,
    \asic/lsdram/msdram/io_dmi_wr_data[152] ,
    \asic/lsdram/msdram/io_dmi_wr_data[151] ,
    \asic/lsdram/msdram/io_dmi_wr_data[150] ,
    \asic/lsdram/msdram/io_dmi_wr_data[149] ,
    \asic/lsdram/msdram/io_dmi_wr_data[148] ,
    \asic/lsdram/msdram/io_dmi_wr_data[147] ,
    \asic/lsdram/msdram/io_dmi_wr_data[146] ,
    \asic/lsdram/msdram/io_dmi_wr_data[145] ,
    \asic/lsdram/msdram/io_dmi_wr_data[144] ,
    \asic/lsdram/msdram/io_dmi_wr_data[143] ,
    \asic/lsdram/msdram/io_dmi_wr_data[142] ,
    \asic/lsdram/msdram/io_dmi_wr_data[141] ,
    \asic/lsdram/msdram/io_dmi_wr_data[140] ,
    \asic/lsdram/msdram/io_dmi_wr_data[139] ,
    \asic/lsdram/msdram/io_dmi_wr_data[138] ,
    \asic/lsdram/msdram/io_dmi_wr_data[137] ,
    \asic/lsdram/msdram/io_dmi_wr_data[136] ,
    \asic/lsdram/msdram/io_dmi_wr_data[135] ,
    \asic/lsdram/msdram/io_dmi_wr_data[134] ,
    \asic/lsdram/msdram/io_dmi_wr_data[133] ,
    \asic/lsdram/msdram/io_dmi_wr_data[132] ,
    \asic/lsdram/msdram/io_dmi_wr_data[131] ,
    \asic/lsdram/msdram/io_dmi_wr_data[130] ,
    \asic/lsdram/msdram/io_dmi_wr_data[129] ,
    \asic/lsdram/msdram/io_dmi_wr_data[128] ,
    \asic/lsdram/msdram/io_dmi_wr_data[127] ,
    \asic/lsdram/msdram/io_dmi_wr_data[126] ,
    \asic/lsdram/msdram/io_dmi_wr_data[125] ,
    \asic/lsdram/msdram/io_dmi_wr_data[124] ,
    \asic/lsdram/msdram/io_dmi_wr_data[123] ,
    \asic/lsdram/msdram/io_dmi_wr_data[122] ,
    \asic/lsdram/msdram/io_dmi_wr_data[121] ,
    \asic/lsdram/msdram/io_dmi_wr_data[120] ,
    \asic/lsdram/msdram/io_dmi_wr_data[119] ,
    \asic/lsdram/msdram/io_dmi_wr_data[118] ,
    \asic/lsdram/msdram/io_dmi_wr_data[117] ,
    \asic/lsdram/msdram/io_dmi_wr_data[116] ,
    \asic/lsdram/msdram/io_dmi_wr_data[115] ,
    \asic/lsdram/msdram/io_dmi_wr_data[114] ,
    \asic/lsdram/msdram/io_dmi_wr_data[113] ,
    \asic/lsdram/msdram/io_dmi_wr_data[112] ,
    \asic/lsdram/msdram/io_dmi_wr_data[111] ,
    \asic/lsdram/msdram/io_dmi_wr_data[110] ,
    \asic/lsdram/msdram/io_dmi_wr_data[109] ,
    \asic/lsdram/msdram/io_dmi_wr_data[108] ,
    \asic/lsdram/msdram/io_dmi_wr_data[107] ,
    \asic/lsdram/msdram/io_dmi_wr_data[106] ,
    \asic/lsdram/msdram/io_dmi_wr_data[105] ,
    \asic/lsdram/msdram/io_dmi_wr_data[104] ,
    \asic/lsdram/msdram/io_dmi_wr_data[103] ,
    \asic/lsdram/msdram/io_dmi_wr_data[102] ,
    \asic/lsdram/msdram/io_dmi_wr_data[101] ,
    \asic/lsdram/msdram/io_dmi_wr_data[100] ,
    \asic/lsdram/msdram/io_dmi_wr_data[99] ,
    \asic/lsdram/msdram/io_dmi_wr_data[98] ,
    \asic/lsdram/msdram/io_dmi_wr_data[97] ,
    \asic/lsdram/msdram/io_dmi_wr_data[96] ,
    \asic/lsdram/msdram/io_dmi_wr_data[95] ,
    \asic/lsdram/msdram/io_dmi_wr_data[94] ,
    \asic/lsdram/msdram/io_dmi_wr_data[93] ,
    \asic/lsdram/msdram/io_dmi_wr_data[92] ,
    \asic/lsdram/msdram/io_dmi_wr_data[91] ,
    \asic/lsdram/msdram/io_dmi_wr_data[90] ,
    \asic/lsdram/msdram/io_dmi_wr_data[89] ,
    \asic/lsdram/msdram/io_dmi_wr_data[88] ,
    \asic/lsdram/msdram/io_dmi_wr_data[87] ,
    \asic/lsdram/msdram/io_dmi_wr_data[86] ,
    \asic/lsdram/msdram/io_dmi_wr_data[85] ,
    \asic/lsdram/msdram/io_dmi_wr_data[84] ,
    \asic/lsdram/msdram/io_dmi_wr_data[83] ,
    \asic/lsdram/msdram/io_dmi_wr_data[82] ,
    \asic/lsdram/msdram/io_dmi_wr_data[81] ,
    \asic/lsdram/msdram/io_dmi_wr_data[80] ,
    \asic/lsdram/msdram/io_dmi_wr_data[79] ,
    \asic/lsdram/msdram/io_dmi_wr_data[78] ,
    \asic/lsdram/msdram/io_dmi_wr_data[77] ,
    \asic/lsdram/msdram/io_dmi_wr_data[76] ,
    \asic/lsdram/msdram/io_dmi_wr_data[75] ,
    \asic/lsdram/msdram/io_dmi_wr_data[74] ,
    \asic/lsdram/msdram/io_dmi_wr_data[73] ,
    \asic/lsdram/msdram/io_dmi_wr_data[72] ,
    \asic/lsdram/msdram/io_dmi_wr_data[71] ,
    \asic/lsdram/msdram/io_dmi_wr_data[70] ,
    \asic/lsdram/msdram/io_dmi_wr_data[69] ,
    \asic/lsdram/msdram/io_dmi_wr_data[68] ,
    \asic/lsdram/msdram/io_dmi_wr_data[67] ,
    \asic/lsdram/msdram/io_dmi_wr_data[66] ,
    \asic/lsdram/msdram/io_dmi_wr_data[65] ,
    \asic/lsdram/msdram/io_dmi_wr_data[64] ,
    \asic/lsdram/msdram/io_dmi_wr_data[63] ,
    \asic/lsdram/msdram/io_dmi_wr_data[62] ,
    \asic/lsdram/msdram/io_dmi_wr_data[61] ,
    \asic/lsdram/msdram/io_dmi_wr_data[60] ,
    \asic/lsdram/msdram/io_dmi_wr_data[59] ,
    \asic/lsdram/msdram/io_dmi_wr_data[58] ,
    \asic/lsdram/msdram/io_dmi_wr_data[57] ,
    \asic/lsdram/msdram/io_dmi_wr_data[56] ,
    \asic/lsdram/msdram/io_dmi_wr_data[55] ,
    \asic/lsdram/msdram/io_dmi_wr_data[54] ,
    \asic/lsdram/msdram/io_dmi_wr_data[53] ,
    \asic/lsdram/msdram/io_dmi_wr_data[52] ,
    \asic/lsdram/msdram/io_dmi_wr_data[51] ,
    \asic/lsdram/msdram/io_dmi_wr_data[50] ,
    \asic/lsdram/msdram/io_dmi_wr_data[49] ,
    \asic/lsdram/msdram/io_dmi_wr_data[48] ,
    \asic/lsdram/msdram/io_dmi_wr_data[47] ,
    \asic/lsdram/msdram/io_dmi_wr_data[46] ,
    \asic/lsdram/msdram/io_dmi_wr_data[45] ,
    \asic/lsdram/msdram/io_dmi_wr_data[44] ,
    \asic/lsdram/msdram/io_dmi_wr_data[43] ,
    \asic/lsdram/msdram/io_dmi_wr_data[42] ,
    \asic/lsdram/msdram/io_dmi_wr_data[41] ,
    \asic/lsdram/msdram/io_dmi_wr_data[40] ,
    \asic/lsdram/msdram/io_dmi_wr_data[39] ,
    \asic/lsdram/msdram/io_dmi_wr_data[38] ,
    \asic/lsdram/msdram/io_dmi_wr_data[37] ,
    \asic/lsdram/msdram/io_dmi_wr_data[36] ,
    \asic/lsdram/msdram/io_dmi_wr_data[35] ,
    \asic/lsdram/msdram/io_dmi_wr_data[34] ,
    \asic/lsdram/msdram/io_dmi_wr_data[33] ,
    \asic/lsdram/msdram/io_dmi_wr_data[32] ,
    \asic/lsdram/msdram/io_dmi_wr_data[31] ,
    \asic/lsdram/msdram/io_dmi_wr_data[30] ,
    \asic/lsdram/msdram/io_dmi_wr_data[29] ,
    \asic/lsdram/msdram/io_dmi_wr_data[28] ,
    \asic/lsdram/msdram/io_dmi_wr_data[27] ,
    \asic/lsdram/msdram/io_dmi_wr_data[26] ,
    \asic/lsdram/msdram/io_dmi_wr_data[25] ,
    \asic/lsdram/msdram/io_dmi_wr_data[24] ,
    \asic/lsdram/msdram/io_dmi_wr_data[23] ,
    \asic/lsdram/msdram/io_dmi_wr_data[22] ,
    \asic/lsdram/msdram/io_dmi_wr_data[21] ,
    \asic/lsdram/msdram/io_dmi_wr_data[20] ,
    \asic/lsdram/msdram/io_dmi_wr_data[19] ,
    \asic/lsdram/msdram/io_dmi_wr_data[18] ,
    \asic/lsdram/msdram/io_dmi_wr_data[17] ,
    \asic/lsdram/msdram/io_dmi_wr_data[16] ,
    \asic/lsdram/msdram/io_dmi_wr_data[15] ,
    \asic/lsdram/msdram/io_dmi_wr_data[14] ,
    \asic/lsdram/msdram/io_dmi_wr_data[13] ,
    \asic/lsdram/msdram/io_dmi_wr_data[12] ,
    \asic/lsdram/msdram/io_dmi_wr_data[11] ,
    \asic/lsdram/msdram/io_dmi_wr_data[10] ,
    \asic/lsdram/msdram/io_dmi_wr_data[9] ,
    \asic/lsdram/msdram/io_dmi_wr_data[8] ,
    \asic/lsdram/msdram/io_dmi_wr_data[7] ,
    \asic/lsdram/msdram/io_dmi_wr_data[6] ,
    \asic/lsdram/msdram/io_dmi_wr_data[5] ,
    \asic/lsdram/msdram/io_dmi_wr_data[4] ,
    \asic/lsdram/msdram/io_dmi_wr_data[3] ,
    \asic/lsdram/msdram/io_dmi_wr_data[2] ,
    \asic/lsdram/msdram/io_dmi_wr_data[1] ,
    \asic/lsdram/msdram/io_dmi_wr_data[0] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[31] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[30] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[29] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[28] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[27] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[26] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[25] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[24] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[23] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[22] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[21] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[20] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[19] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[18] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[17] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[16] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[15] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[14] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[13] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[12] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[11] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[10] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[9] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[8] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[7] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[6] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[5] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[4] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[3] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[2] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[1] ,
    \asic/lsdram/msdram/io_dmi_wr_data_mask[0] ,
    \asic/lsdram/msdram/io_dmi_rd_data[255] ,
    \asic/lsdram/msdram/io_dmi_rd_data[254] ,
    \asic/lsdram/msdram/io_dmi_rd_data[253] ,
    \asic/lsdram/msdram/io_dmi_rd_data[252] ,
    \asic/lsdram/msdram/io_dmi_rd_data[251] ,
    \asic/lsdram/msdram/io_dmi_rd_data[250] ,
    \asic/lsdram/msdram/io_dmi_rd_data[249] ,
    \asic/lsdram/msdram/io_dmi_rd_data[248] ,
    \asic/lsdram/msdram/io_dmi_rd_data[247] ,
    \asic/lsdram/msdram/io_dmi_rd_data[246] ,
    \asic/lsdram/msdram/io_dmi_rd_data[245] ,
    \asic/lsdram/msdram/io_dmi_rd_data[244] ,
    \asic/lsdram/msdram/io_dmi_rd_data[243] ,
    \asic/lsdram/msdram/io_dmi_rd_data[242] ,
    \asic/lsdram/msdram/io_dmi_rd_data[241] ,
    \asic/lsdram/msdram/io_dmi_rd_data[240] ,
    \asic/lsdram/msdram/io_dmi_rd_data[239] ,
    \asic/lsdram/msdram/io_dmi_rd_data[238] ,
    \asic/lsdram/msdram/io_dmi_rd_data[237] ,
    \asic/lsdram/msdram/io_dmi_rd_data[236] ,
    \asic/lsdram/msdram/io_dmi_rd_data[235] ,
    \asic/lsdram/msdram/io_dmi_rd_data[234] ,
    \asic/lsdram/msdram/io_dmi_rd_data[233] ,
    \asic/lsdram/msdram/io_dmi_rd_data[232] ,
    \asic/lsdram/msdram/io_dmi_rd_data[231] ,
    \asic/lsdram/msdram/io_dmi_rd_data[230] ,
    \asic/lsdram/msdram/io_dmi_rd_data[229] ,
    \asic/lsdram/msdram/io_dmi_rd_data[228] ,
    \asic/lsdram/msdram/io_dmi_rd_data[227] ,
    \asic/lsdram/msdram/io_dmi_rd_data[226] ,
    \asic/lsdram/msdram/io_dmi_rd_data[225] ,
    \asic/lsdram/msdram/io_dmi_rd_data[224] ,
    \asic/lsdram/msdram/io_dmi_rd_data[223] ,
    \asic/lsdram/msdram/io_dmi_rd_data[222] ,
    \asic/lsdram/msdram/io_dmi_rd_data[221] ,
    \asic/lsdram/msdram/io_dmi_rd_data[220] ,
    \asic/lsdram/msdram/io_dmi_rd_data[219] ,
    \asic/lsdram/msdram/io_dmi_rd_data[218] ,
    \asic/lsdram/msdram/io_dmi_rd_data[217] ,
    \asic/lsdram/msdram/io_dmi_rd_data[216] ,
    \asic/lsdram/msdram/io_dmi_rd_data[215] ,
    \asic/lsdram/msdram/io_dmi_rd_data[214] ,
    \asic/lsdram/msdram/io_dmi_rd_data[213] ,
    \asic/lsdram/msdram/io_dmi_rd_data[212] ,
    \asic/lsdram/msdram/io_dmi_rd_data[211] ,
    \asic/lsdram/msdram/io_dmi_rd_data[210] ,
    \asic/lsdram/msdram/io_dmi_rd_data[209] ,
    \asic/lsdram/msdram/io_dmi_rd_data[208] ,
    \asic/lsdram/msdram/io_dmi_rd_data[207] ,
    \asic/lsdram/msdram/io_dmi_rd_data[206] ,
    \asic/lsdram/msdram/io_dmi_rd_data[205] ,
    \asic/lsdram/msdram/io_dmi_rd_data[204] ,
    \asic/lsdram/msdram/io_dmi_rd_data[203] ,
    \asic/lsdram/msdram/io_dmi_rd_data[202] ,
    \asic/lsdram/msdram/io_dmi_rd_data[201] ,
    \asic/lsdram/msdram/io_dmi_rd_data[200] ,
    \asic/lsdram/msdram/io_dmi_rd_data[199] ,
    \asic/lsdram/msdram/io_dmi_rd_data[198] ,
    \asic/lsdram/msdram/io_dmi_rd_data[197] ,
    \asic/lsdram/msdram/io_dmi_rd_data[196] ,
    \asic/lsdram/msdram/io_dmi_rd_data[195] ,
    \asic/lsdram/msdram/io_dmi_rd_data[194] ,
    \asic/lsdram/msdram/io_dmi_rd_data[193] ,
    \asic/lsdram/msdram/io_dmi_rd_data[192] ,
    \asic/lsdram/msdram/io_dmi_rd_data[191] ,
    \asic/lsdram/msdram/io_dmi_rd_data[190] ,
    \asic/lsdram/msdram/io_dmi_rd_data[189] ,
    \asic/lsdram/msdram/io_dmi_rd_data[188] ,
    \asic/lsdram/msdram/io_dmi_rd_data[187] ,
    \asic/lsdram/msdram/io_dmi_rd_data[186] ,
    \asic/lsdram/msdram/io_dmi_rd_data[185] ,
    \asic/lsdram/msdram/io_dmi_rd_data[184] ,
    \asic/lsdram/msdram/io_dmi_rd_data[183] ,
    \asic/lsdram/msdram/io_dmi_rd_data[182] ,
    \asic/lsdram/msdram/io_dmi_rd_data[181] ,
    \asic/lsdram/msdram/io_dmi_rd_data[180] ,
    \asic/lsdram/msdram/io_dmi_rd_data[179] ,
    \asic/lsdram/msdram/io_dmi_rd_data[178] ,
    \asic/lsdram/msdram/io_dmi_rd_data[177] ,
    \asic/lsdram/msdram/io_dmi_rd_data[176] ,
    \asic/lsdram/msdram/io_dmi_rd_data[175] ,
    \asic/lsdram/msdram/io_dmi_rd_data[174] ,
    \asic/lsdram/msdram/io_dmi_rd_data[173] ,
    \asic/lsdram/msdram/io_dmi_rd_data[172] ,
    \asic/lsdram/msdram/io_dmi_rd_data[171] ,
    \asic/lsdram/msdram/io_dmi_rd_data[170] ,
    \asic/lsdram/msdram/io_dmi_rd_data[169] ,
    \asic/lsdram/msdram/io_dmi_rd_data[168] ,
    \asic/lsdram/msdram/io_dmi_rd_data[167] ,
    \asic/lsdram/msdram/io_dmi_rd_data[166] ,
    \asic/lsdram/msdram/io_dmi_rd_data[165] ,
    \asic/lsdram/msdram/io_dmi_rd_data[164] ,
    \asic/lsdram/msdram/io_dmi_rd_data[163] ,
    \asic/lsdram/msdram/io_dmi_rd_data[162] ,
    \asic/lsdram/msdram/io_dmi_rd_data[161] ,
    \asic/lsdram/msdram/io_dmi_rd_data[160] ,
    \asic/lsdram/msdram/io_dmi_rd_data[159] ,
    \asic/lsdram/msdram/io_dmi_rd_data[158] ,
    \asic/lsdram/msdram/io_dmi_rd_data[157] ,
    \asic/lsdram/msdram/io_dmi_rd_data[156] ,
    \asic/lsdram/msdram/io_dmi_rd_data[155] ,
    \asic/lsdram/msdram/io_dmi_rd_data[154] ,
    \asic/lsdram/msdram/io_dmi_rd_data[153] ,
    \asic/lsdram/msdram/io_dmi_rd_data[152] ,
    \asic/lsdram/msdram/io_dmi_rd_data[151] ,
    \asic/lsdram/msdram/io_dmi_rd_data[150] ,
    \asic/lsdram/msdram/io_dmi_rd_data[149] ,
    \asic/lsdram/msdram/io_dmi_rd_data[148] ,
    \asic/lsdram/msdram/io_dmi_rd_data[147] ,
    \asic/lsdram/msdram/io_dmi_rd_data[146] ,
    \asic/lsdram/msdram/io_dmi_rd_data[145] ,
    \asic/lsdram/msdram/io_dmi_rd_data[144] ,
    \asic/lsdram/msdram/io_dmi_rd_data[143] ,
    \asic/lsdram/msdram/io_dmi_rd_data[142] ,
    \asic/lsdram/msdram/io_dmi_rd_data[141] ,
    \asic/lsdram/msdram/io_dmi_rd_data[140] ,
    \asic/lsdram/msdram/io_dmi_rd_data[139] ,
    \asic/lsdram/msdram/io_dmi_rd_data[138] ,
    \asic/lsdram/msdram/io_dmi_rd_data[137] ,
    \asic/lsdram/msdram/io_dmi_rd_data[136] ,
    \asic/lsdram/msdram/io_dmi_rd_data[135] ,
    \asic/lsdram/msdram/io_dmi_rd_data[134] ,
    \asic/lsdram/msdram/io_dmi_rd_data[133] ,
    \asic/lsdram/msdram/io_dmi_rd_data[132] ,
    \asic/lsdram/msdram/io_dmi_rd_data[131] ,
    \asic/lsdram/msdram/io_dmi_rd_data[130] ,
    \asic/lsdram/msdram/io_dmi_rd_data[129] ,
    \asic/lsdram/msdram/io_dmi_rd_data[128] ,
    \asic/lsdram/msdram/io_dmi_rd_data[127] ,
    \asic/lsdram/msdram/io_dmi_rd_data[126] ,
    \asic/lsdram/msdram/io_dmi_rd_data[125] ,
    \asic/lsdram/msdram/io_dmi_rd_data[124] ,
    \asic/lsdram/msdram/io_dmi_rd_data[123] ,
    \asic/lsdram/msdram/io_dmi_rd_data[122] ,
    \asic/lsdram/msdram/io_dmi_rd_data[121] ,
    \asic/lsdram/msdram/io_dmi_rd_data[120] ,
    \asic/lsdram/msdram/io_dmi_rd_data[119] ,
    \asic/lsdram/msdram/io_dmi_rd_data[118] ,
    \asic/lsdram/msdram/io_dmi_rd_data[117] ,
    \asic/lsdram/msdram/io_dmi_rd_data[116] ,
    \asic/lsdram/msdram/io_dmi_rd_data[115] ,
    \asic/lsdram/msdram/io_dmi_rd_data[114] ,
    \asic/lsdram/msdram/io_dmi_rd_data[113] ,
    \asic/lsdram/msdram/io_dmi_rd_data[112] ,
    \asic/lsdram/msdram/io_dmi_rd_data[111] ,
    \asic/lsdram/msdram/io_dmi_rd_data[110] ,
    \asic/lsdram/msdram/io_dmi_rd_data[109] ,
    \asic/lsdram/msdram/io_dmi_rd_data[108] ,
    \asic/lsdram/msdram/io_dmi_rd_data[107] ,
    \asic/lsdram/msdram/io_dmi_rd_data[106] ,
    \asic/lsdram/msdram/io_dmi_rd_data[105] ,
    \asic/lsdram/msdram/io_dmi_rd_data[104] ,
    \asic/lsdram/msdram/io_dmi_rd_data[103] ,
    \asic/lsdram/msdram/io_dmi_rd_data[102] ,
    \asic/lsdram/msdram/io_dmi_rd_data[101] ,
    \asic/lsdram/msdram/io_dmi_rd_data[100] ,
    \asic/lsdram/msdram/io_dmi_rd_data[99] ,
    \asic/lsdram/msdram/io_dmi_rd_data[98] ,
    \asic/lsdram/msdram/io_dmi_rd_data[97] ,
    \asic/lsdram/msdram/io_dmi_rd_data[96] ,
    \asic/lsdram/msdram/io_dmi_rd_data[95] ,
    \asic/lsdram/msdram/io_dmi_rd_data[94] ,
    \asic/lsdram/msdram/io_dmi_rd_data[93] ,
    \asic/lsdram/msdram/io_dmi_rd_data[92] ,
    \asic/lsdram/msdram/io_dmi_rd_data[91] ,
    \asic/lsdram/msdram/io_dmi_rd_data[90] ,
    \asic/lsdram/msdram/io_dmi_rd_data[89] ,
    \asic/lsdram/msdram/io_dmi_rd_data[88] ,
    \asic/lsdram/msdram/io_dmi_rd_data[87] ,
    \asic/lsdram/msdram/io_dmi_rd_data[86] ,
    \asic/lsdram/msdram/io_dmi_rd_data[85] ,
    \asic/lsdram/msdram/io_dmi_rd_data[84] ,
    \asic/lsdram/msdram/io_dmi_rd_data[83] ,
    \asic/lsdram/msdram/io_dmi_rd_data[82] ,
    \asic/lsdram/msdram/io_dmi_rd_data[81] ,
    \asic/lsdram/msdram/io_dmi_rd_data[80] ,
    \asic/lsdram/msdram/io_dmi_rd_data[79] ,
    \asic/lsdram/msdram/io_dmi_rd_data[78] ,
    \asic/lsdram/msdram/io_dmi_rd_data[77] ,
    \asic/lsdram/msdram/io_dmi_rd_data[76] ,
    \asic/lsdram/msdram/io_dmi_rd_data[75] ,
    \asic/lsdram/msdram/io_dmi_rd_data[74] ,
    \asic/lsdram/msdram/io_dmi_rd_data[73] ,
    \asic/lsdram/msdram/io_dmi_rd_data[72] ,
    \asic/lsdram/msdram/io_dmi_rd_data[71] ,
    \asic/lsdram/msdram/io_dmi_rd_data[70] ,
    \asic/lsdram/msdram/io_dmi_rd_data[69] ,
    \asic/lsdram/msdram/io_dmi_rd_data[68] ,
    \asic/lsdram/msdram/io_dmi_rd_data[67] ,
    \asic/lsdram/msdram/io_dmi_rd_data[66] ,
    \asic/lsdram/msdram/io_dmi_rd_data[65] ,
    \asic/lsdram/msdram/io_dmi_rd_data[64] ,
    \asic/lsdram/msdram/io_dmi_rd_data[63] ,
    \asic/lsdram/msdram/io_dmi_rd_data[62] ,
    \asic/lsdram/msdram/io_dmi_rd_data[61] ,
    \asic/lsdram/msdram/io_dmi_rd_data[60] ,
    \asic/lsdram/msdram/io_dmi_rd_data[59] ,
    \asic/lsdram/msdram/io_dmi_rd_data[58] ,
    \asic/lsdram/msdram/io_dmi_rd_data[57] ,
    \asic/lsdram/msdram/io_dmi_rd_data[56] ,
    \asic/lsdram/msdram/io_dmi_rd_data[55] ,
    \asic/lsdram/msdram/io_dmi_rd_data[54] ,
    \asic/lsdram/msdram/io_dmi_rd_data[53] ,
    \asic/lsdram/msdram/io_dmi_rd_data[52] ,
    \asic/lsdram/msdram/io_dmi_rd_data[51] ,
    \asic/lsdram/msdram/io_dmi_rd_data[50] ,
    \asic/lsdram/msdram/io_dmi_rd_data[49] ,
    \asic/lsdram/msdram/io_dmi_rd_data[48] ,
    \asic/lsdram/msdram/io_dmi_rd_data[47] ,
    \asic/lsdram/msdram/io_dmi_rd_data[46] ,
    \asic/lsdram/msdram/io_dmi_rd_data[45] ,
    \asic/lsdram/msdram/io_dmi_rd_data[44] ,
    \asic/lsdram/msdram/io_dmi_rd_data[43] ,
    \asic/lsdram/msdram/io_dmi_rd_data[42] ,
    \asic/lsdram/msdram/io_dmi_rd_data[41] ,
    \asic/lsdram/msdram/io_dmi_rd_data[40] ,
    \asic/lsdram/msdram/io_dmi_rd_data[39] ,
    \asic/lsdram/msdram/io_dmi_rd_data[38] ,
    \asic/lsdram/msdram/io_dmi_rd_data[37] ,
    \asic/lsdram/msdram/io_dmi_rd_data[36] ,
    \asic/lsdram/msdram/io_dmi_rd_data[35] ,
    \asic/lsdram/msdram/io_dmi_rd_data[34] ,
    \asic/lsdram/msdram/io_dmi_rd_data[33] ,
    \asic/lsdram/msdram/io_dmi_rd_data[32] ,
    \asic/lsdram/msdram/io_dmi_rd_data[31] ,
    \asic/lsdram/msdram/io_dmi_rd_data[30] ,
    \asic/lsdram/msdram/io_dmi_rd_data[29] ,
    \asic/lsdram/msdram/io_dmi_rd_data[28] ,
    \asic/lsdram/msdram/io_dmi_rd_data[27] ,
    \asic/lsdram/msdram/io_dmi_rd_data[26] ,
    \asic/lsdram/msdram/io_dmi_rd_data[25] ,
    \asic/lsdram/msdram/io_dmi_rd_data[24] ,
    \asic/lsdram/msdram/io_dmi_rd_data[23] ,
    \asic/lsdram/msdram/io_dmi_rd_data[22] ,
    \asic/lsdram/msdram/io_dmi_rd_data[21] ,
    \asic/lsdram/msdram/io_dmi_rd_data[20] ,
    \asic/lsdram/msdram/io_dmi_rd_data[19] ,
    \asic/lsdram/msdram/io_dmi_rd_data[18] ,
    \asic/lsdram/msdram/io_dmi_rd_data[17] ,
    \asic/lsdram/msdram/io_dmi_rd_data[16] ,
    \asic/lsdram/msdram/io_dmi_rd_data[15] ,
    \asic/lsdram/msdram/io_dmi_rd_data[14] ,
    \asic/lsdram/msdram/io_dmi_rd_data[13] ,
    \asic/lsdram/msdram/io_dmi_rd_data[12] ,
    \asic/lsdram/msdram/io_dmi_rd_data[11] ,
    \asic/lsdram/msdram/io_dmi_rd_data[10] ,
    \asic/lsdram/msdram/io_dmi_rd_data[9] ,
    \asic/lsdram/msdram/io_dmi_rd_data[8] ,
    \asic/lsdram/msdram/io_dmi_rd_data[7] ,
    \asic/lsdram/msdram/io_dmi_rd_data[6] ,
    \asic/lsdram/msdram/io_dmi_rd_data[5] ,
    \asic/lsdram/msdram/io_dmi_rd_data[4] ,
    \asic/lsdram/msdram/io_dmi_rd_data[3] ,
    \asic/lsdram/msdram/io_dmi_rd_data[2] ,
    \asic/lsdram/msdram/io_dmi_rd_data[1] ,
    \asic/lsdram/msdram/io_dmi_rd_data[0] ,
    \asic/lsdram/msdram/io_in_rdata_r[255] ,
    \asic/lsdram/msdram/io_in_rdata_r[254] ,
    \asic/lsdram/msdram/io_in_rdata_r[253] ,
    \asic/lsdram/msdram/io_in_rdata_r[252] ,
    \asic/lsdram/msdram/io_in_rdata_r[251] ,
    \asic/lsdram/msdram/io_in_rdata_r[250] ,
    \asic/lsdram/msdram/io_in_rdata_r[249] ,
    \asic/lsdram/msdram/io_in_rdata_r[248] ,
    \asic/lsdram/msdram/io_in_rdata_r[247] ,
    \asic/lsdram/msdram/io_in_rdata_r[246] ,
    \asic/lsdram/msdram/io_in_rdata_r[245] ,
    \asic/lsdram/msdram/io_in_rdata_r[244] ,
    \asic/lsdram/msdram/io_in_rdata_r[243] ,
    \asic/lsdram/msdram/io_in_rdata_r[242] ,
    \asic/lsdram/msdram/io_in_rdata_r[241] ,
    \asic/lsdram/msdram/io_in_rdata_r[240] ,
    \asic/lsdram/msdram/io_in_rdata_r[239] ,
    \asic/lsdram/msdram/io_in_rdata_r[238] ,
    \asic/lsdram/msdram/io_in_rdata_r[237] ,
    \asic/lsdram/msdram/io_in_rdata_r[236] ,
    \asic/lsdram/msdram/io_in_rdata_r[235] ,
    \asic/lsdram/msdram/io_in_rdata_r[234] ,
    \asic/lsdram/msdram/io_in_rdata_r[233] ,
    \asic/lsdram/msdram/io_in_rdata_r[232] ,
    \asic/lsdram/msdram/io_in_rdata_r[231] ,
    \asic/lsdram/msdram/io_in_rdata_r[230] ,
    \asic/lsdram/msdram/io_in_rdata_r[229] ,
    \asic/lsdram/msdram/io_in_rdata_r[228] ,
    \asic/lsdram/msdram/io_in_rdata_r[227] ,
    \asic/lsdram/msdram/io_in_rdata_r[226] ,
    \asic/lsdram/msdram/io_in_rdata_r[225] ,
    \asic/lsdram/msdram/io_in_rdata_r[224] ,
    \asic/lsdram/msdram/io_in_rdata_r[223] ,
    \asic/lsdram/msdram/io_in_rdata_r[222] ,
    \asic/lsdram/msdram/io_in_rdata_r[221] ,
    \asic/lsdram/msdram/io_in_rdata_r[220] ,
    \asic/lsdram/msdram/io_in_rdata_r[219] ,
    \asic/lsdram/msdram/io_in_rdata_r[218] ,
    \asic/lsdram/msdram/io_in_rdata_r[217] ,
    \asic/lsdram/msdram/io_in_rdata_r[216] ,
    \asic/lsdram/msdram/io_in_rdata_r[215] ,
    \asic/lsdram/msdram/io_in_rdata_r[214] ,
    \asic/lsdram/msdram/io_in_rdata_r[213] ,
    \asic/lsdram/msdram/io_in_rdata_r[212] ,
    \asic/lsdram/msdram/io_in_rdata_r[211] ,
    \asic/lsdram/msdram/io_in_rdata_r[210] ,
    \asic/lsdram/msdram/io_in_rdata_r[209] ,
    \asic/lsdram/msdram/io_in_rdata_r[208] ,
    \asic/lsdram/msdram/io_in_rdata_r[207] ,
    \asic/lsdram/msdram/io_in_rdata_r[206] ,
    \asic/lsdram/msdram/io_in_rdata_r[205] ,
    \asic/lsdram/msdram/io_in_rdata_r[204] ,
    \asic/lsdram/msdram/io_in_rdata_r[203] ,
    \asic/lsdram/msdram/io_in_rdata_r[202] ,
    \asic/lsdram/msdram/io_in_rdata_r[201] ,
    \asic/lsdram/msdram/io_in_rdata_r[200] ,
    \asic/lsdram/msdram/io_in_rdata_r[199] ,
    \asic/lsdram/msdram/io_in_rdata_r[198] ,
    \asic/lsdram/msdram/io_in_rdata_r[197] ,
    \asic/lsdram/msdram/io_in_rdata_r[196] ,
    \asic/lsdram/msdram/io_in_rdata_r[195] ,
    \asic/lsdram/msdram/io_in_rdata_r[194] ,
    \asic/lsdram/msdram/io_in_rdata_r[193] ,
    \asic/lsdram/msdram/io_in_rdata_r[192] ,
    \asic/lsdram/msdram/io_in_rdata_r[191] ,
    \asic/lsdram/msdram/io_in_rdata_r[190] ,
    \asic/lsdram/msdram/io_in_rdata_r[189] ,
    \asic/lsdram/msdram/io_in_rdata_r[188] ,
    \asic/lsdram/msdram/io_in_rdata_r[187] ,
    \asic/lsdram/msdram/io_in_rdata_r[186] ,
    \asic/lsdram/msdram/io_in_rdata_r[185] ,
    \asic/lsdram/msdram/io_in_rdata_r[184] ,
    \asic/lsdram/msdram/io_in_rdata_r[183] ,
    \asic/lsdram/msdram/io_in_rdata_r[182] ,
    \asic/lsdram/msdram/io_in_rdata_r[181] ,
    \asic/lsdram/msdram/io_in_rdata_r[180] ,
    \asic/lsdram/msdram/io_in_rdata_r[179] ,
    \asic/lsdram/msdram/io_in_rdata_r[178] ,
    \asic/lsdram/msdram/io_in_rdata_r[177] ,
    \asic/lsdram/msdram/io_in_rdata_r[176] ,
    \asic/lsdram/msdram/io_in_rdata_r[175] ,
    \asic/lsdram/msdram/io_in_rdata_r[174] ,
    \asic/lsdram/msdram/io_in_rdata_r[173] ,
    \asic/lsdram/msdram/io_in_rdata_r[172] ,
    \asic/lsdram/msdram/io_in_rdata_r[171] ,
    \asic/lsdram/msdram/io_in_rdata_r[170] ,
    \asic/lsdram/msdram/io_in_rdata_r[169] ,
    \asic/lsdram/msdram/io_in_rdata_r[168] ,
    \asic/lsdram/msdram/io_in_rdata_r[167] ,
    \asic/lsdram/msdram/io_in_rdata_r[166] ,
    \asic/lsdram/msdram/io_in_rdata_r[165] ,
    \asic/lsdram/msdram/io_in_rdata_r[164] ,
    \asic/lsdram/msdram/io_in_rdata_r[163] ,
    \asic/lsdram/msdram/io_in_rdata_r[162] ,
    \asic/lsdram/msdram/io_in_rdata_r[161] ,
    \asic/lsdram/msdram/io_in_rdata_r[160] ,
    \asic/lsdram/msdram/io_in_rdata_r[159] ,
    \asic/lsdram/msdram/io_in_rdata_r[158] ,
    \asic/lsdram/msdram/io_in_rdata_r[157] ,
    \asic/lsdram/msdram/io_in_rdata_r[156] ,
    \asic/lsdram/msdram/io_in_rdata_r[155] ,
    \asic/lsdram/msdram/io_in_rdata_r[154] ,
    \asic/lsdram/msdram/io_in_rdata_r[153] ,
    \asic/lsdram/msdram/io_in_rdata_r[152] ,
    \asic/lsdram/msdram/io_in_rdata_r[151] ,
    \asic/lsdram/msdram/io_in_rdata_r[150] ,
    \asic/lsdram/msdram/io_in_rdata_r[149] ,
    \asic/lsdram/msdram/io_in_rdata_r[148] ,
    \asic/lsdram/msdram/io_in_rdata_r[147] ,
    \asic/lsdram/msdram/io_in_rdata_r[146] ,
    \asic/lsdram/msdram/io_in_rdata_r[145] ,
    \asic/lsdram/msdram/io_in_rdata_r[144] ,
    \asic/lsdram/msdram/io_in_rdata_r[143] ,
    \asic/lsdram/msdram/io_in_rdata_r[142] ,
    \asic/lsdram/msdram/io_in_rdata_r[141] ,
    \asic/lsdram/msdram/io_in_rdata_r[140] ,
    \asic/lsdram/msdram/io_in_rdata_r[139] ,
    \asic/lsdram/msdram/io_in_rdata_r[138] ,
    \asic/lsdram/msdram/io_in_rdata_r[137] ,
    \asic/lsdram/msdram/io_in_rdata_r[136] ,
    \asic/lsdram/msdram/io_in_rdata_r[135] ,
    \asic/lsdram/msdram/io_in_rdata_r[134] ,
    \asic/lsdram/msdram/io_in_rdata_r[133] ,
    \asic/lsdram/msdram/io_in_rdata_r[132] ,
    \asic/lsdram/msdram/io_in_rdata_r[131] ,
    \asic/lsdram/msdram/io_in_rdata_r[130] ,
    \asic/lsdram/msdram/io_in_rdata_r[129] ,
    \asic/lsdram/msdram/io_in_rdata_r[128] ,
    \asic/lsdram/msdram/io_in_rdata_r[127] ,
    \asic/lsdram/msdram/io_in_rdata_r[126] ,
    \asic/lsdram/msdram/io_in_rdata_r[125] ,
    \asic/lsdram/msdram/io_in_rdata_r[124] ,
    \asic/lsdram/msdram/io_in_rdata_r[123] ,
    \asic/lsdram/msdram/io_in_rdata_r[122] ,
    \asic/lsdram/msdram/io_in_rdata_r[121] ,
    \asic/lsdram/msdram/io_in_rdata_r[120] ,
    \asic/lsdram/msdram/io_in_rdata_r[119] ,
    \asic/lsdram/msdram/io_in_rdata_r[118] ,
    \asic/lsdram/msdram/io_in_rdata_r[117] ,
    \asic/lsdram/msdram/io_in_rdata_r[116] ,
    \asic/lsdram/msdram/io_in_rdata_r[115] ,
    \asic/lsdram/msdram/io_in_rdata_r[114] ,
    \asic/lsdram/msdram/io_in_rdata_r[113] ,
    \asic/lsdram/msdram/io_in_rdata_r[112] ,
    \asic/lsdram/msdram/io_in_rdata_r[111] ,
    \asic/lsdram/msdram/io_in_rdata_r[110] ,
    \asic/lsdram/msdram/io_in_rdata_r[109] ,
    \asic/lsdram/msdram/io_in_rdata_r[108] ,
    \asic/lsdram/msdram/io_in_rdata_r[107] ,
    \asic/lsdram/msdram/io_in_rdata_r[106] ,
    \asic/lsdram/msdram/io_in_rdata_r[105] ,
    \asic/lsdram/msdram/io_in_rdata_r[104] ,
    \asic/lsdram/msdram/io_in_rdata_r[103] ,
    \asic/lsdram/msdram/io_in_rdata_r[102] ,
    \asic/lsdram/msdram/io_in_rdata_r[101] ,
    \asic/lsdram/msdram/io_in_rdata_r[100] ,
    \asic/lsdram/msdram/io_in_rdata_r[99] ,
    \asic/lsdram/msdram/io_in_rdata_r[98] ,
    \asic/lsdram/msdram/io_in_rdata_r[97] ,
    \asic/lsdram/msdram/io_in_rdata_r[96] ,
    \asic/lsdram/msdram/io_in_rdata_r[95] ,
    \asic/lsdram/msdram/io_in_rdata_r[94] ,
    \asic/lsdram/msdram/io_in_rdata_r[93] ,
    \asic/lsdram/msdram/io_in_rdata_r[92] ,
    \asic/lsdram/msdram/io_in_rdata_r[91] ,
    \asic/lsdram/msdram/io_in_rdata_r[90] ,
    \asic/lsdram/msdram/io_in_rdata_r[89] ,
    \asic/lsdram/msdram/io_in_rdata_r[88] ,
    \asic/lsdram/msdram/io_in_rdata_r[87] ,
    \asic/lsdram/msdram/io_in_rdata_r[86] ,
    \asic/lsdram/msdram/io_in_rdata_r[85] ,
    \asic/lsdram/msdram/io_in_rdata_r[84] ,
    \asic/lsdram/msdram/io_in_rdata_r[83] ,
    \asic/lsdram/msdram/io_in_rdata_r[82] ,
    \asic/lsdram/msdram/io_in_rdata_r[81] ,
    \asic/lsdram/msdram/io_in_rdata_r[80] ,
    \asic/lsdram/msdram/io_in_rdata_r[79] ,
    \asic/lsdram/msdram/io_in_rdata_r[78] ,
    \asic/lsdram/msdram/io_in_rdata_r[77] ,
    \asic/lsdram/msdram/io_in_rdata_r[76] ,
    \asic/lsdram/msdram/io_in_rdata_r[75] ,
    \asic/lsdram/msdram/io_in_rdata_r[74] ,
    \asic/lsdram/msdram/io_in_rdata_r[73] ,
    \asic/lsdram/msdram/io_in_rdata_r[72] ,
    \asic/lsdram/msdram/io_in_rdata_r[71] ,
    \asic/lsdram/msdram/io_in_rdata_r[70] ,
    \asic/lsdram/msdram/io_in_rdata_r[69] ,
    \asic/lsdram/msdram/io_in_rdata_r[68] ,
    \asic/lsdram/msdram/io_in_rdata_r[67] ,
    \asic/lsdram/msdram/io_in_rdata_r[66] ,
    \asic/lsdram/msdram/io_in_rdata_r[65] ,
    \asic/lsdram/msdram/io_in_rdata_r[64] ,
    \asic/lsdram/msdram/io_in_rdata_r[63] ,
    \asic/lsdram/msdram/io_in_rdata_r[62] ,
    \asic/lsdram/msdram/io_in_rdata_r[61] ,
    \asic/lsdram/msdram/io_in_rdata_r[60] ,
    \asic/lsdram/msdram/io_in_rdata_r[59] ,
    \asic/lsdram/msdram/io_in_rdata_r[58] ,
    \asic/lsdram/msdram/io_in_rdata_r[57] ,
    \asic/lsdram/msdram/io_in_rdata_r[56] ,
    \asic/lsdram/msdram/io_in_rdata_r[55] ,
    \asic/lsdram/msdram/io_in_rdata_r[54] ,
    \asic/lsdram/msdram/io_in_rdata_r[53] ,
    \asic/lsdram/msdram/io_in_rdata_r[52] ,
    \asic/lsdram/msdram/io_in_rdata_r[51] ,
    \asic/lsdram/msdram/io_in_rdata_r[50] ,
    \asic/lsdram/msdram/io_in_rdata_r[49] ,
    \asic/lsdram/msdram/io_in_rdata_r[48] ,
    \asic/lsdram/msdram/io_in_rdata_r[47] ,
    \asic/lsdram/msdram/io_in_rdata_r[46] ,
    \asic/lsdram/msdram/io_in_rdata_r[45] ,
    \asic/lsdram/msdram/io_in_rdata_r[44] ,
    \asic/lsdram/msdram/io_in_rdata_r[43] ,
    \asic/lsdram/msdram/io_in_rdata_r[42] ,
    \asic/lsdram/msdram/io_in_rdata_r[41] ,
    \asic/lsdram/msdram/io_in_rdata_r[40] ,
    \asic/lsdram/msdram/io_in_rdata_r[39] ,
    \asic/lsdram/msdram/io_in_rdata_r[38] ,
    \asic/lsdram/msdram/io_in_rdata_r[37] ,
    \asic/lsdram/msdram/io_in_rdata_r[36] ,
    \asic/lsdram/msdram/io_in_rdata_r[35] ,
    \asic/lsdram/msdram/io_in_rdata_r[34] ,
    \asic/lsdram/msdram/io_in_rdata_r[33] ,
    \asic/lsdram/msdram/io_in_rdata_r[32] ,
    \asic/lsdram/msdram/io_in_rdata_r[31] ,
    \asic/lsdram/msdram/io_in_rdata_r[30] ,
    \asic/lsdram/msdram/io_in_rdata_r[29] ,
    \asic/lsdram/msdram/io_in_rdata_r[28] ,
    \asic/lsdram/msdram/io_in_rdata_r[27] ,
    \asic/lsdram/msdram/io_in_rdata_r[26] ,
    \asic/lsdram/msdram/io_in_rdata_r[25] ,
    \asic/lsdram/msdram/io_in_rdata_r[24] ,
    \asic/lsdram/msdram/io_in_rdata_r[23] ,
    \asic/lsdram/msdram/io_in_rdata_r[22] ,
    \asic/lsdram/msdram/io_in_rdata_r[21] ,
    \asic/lsdram/msdram/io_in_rdata_r[20] ,
    \asic/lsdram/msdram/io_in_rdata_r[19] ,
    \asic/lsdram/msdram/io_in_rdata_r[18] ,
    \asic/lsdram/msdram/io_in_rdata_r[17] ,
    \asic/lsdram/msdram/io_in_rdata_r[16] ,
    \asic/lsdram/msdram/io_in_rdata_r[15] ,
    \asic/lsdram/msdram/io_in_rdata_r[14] ,
    \asic/lsdram/msdram/io_in_rdata_r[13] ,
    \asic/lsdram/msdram/io_in_rdata_r[12] ,
    \asic/lsdram/msdram/io_in_rdata_r[11] ,
    \asic/lsdram/msdram/io_in_rdata_r[10] ,
    \asic/lsdram/msdram/io_in_rdata_r[9] ,
    \asic/lsdram/msdram/io_in_rdata_r[8] ,
    \asic/lsdram/msdram/io_in_rdata_r[7] ,
    \asic/lsdram/msdram/io_in_rdata_r[6] ,
    \asic/lsdram/msdram/io_in_rdata_r[5] ,
    \asic/lsdram/msdram/io_in_rdata_r[4] ,
    \asic/lsdram/msdram/io_in_rdata_r[3] ,
    \asic/lsdram/msdram/io_in_rdata_r[2] ,
    \asic/lsdram/msdram/io_in_rdata_r[1] ,
    \asic/lsdram/msdram/io_in_rdata_r[0] ,
    \asic/lsdram/msdram/io_clk_out ,
    \asic/lsdram/msdram/io_in_awready ,
    \asic/lsdram/msdram/io_in_awvalid ,
    \asic/lsdram/msdram/io_in_wready ,
    \asic/lsdram/msdram/io_in_wvalid ,
    \asic/lsdram/msdram/io_in_bready ,
    \asic/lsdram/msdram/io_in_bvalid ,
    \asic/lsdram/msdram/io_in_arready ,
    \asic/lsdram/msdram/io_in_arvalid ,
    \asic/lsdram/msdram/io_in_rready ,
    \asic/lsdram/msdram/io_in_rvalid ,
    \asic/lsdram/msdram/io_dmi_cmd_en ,
    \asic/lsdram/msdram/io_dmi_wr_data_en ,
    \asic/lsdram/msdram/io_dmi_wr_data_end ,
    \asic/lsdram/msdram/io_dmi_clk_out ,
    \asic/lsdram/msdram/io_dmi_init_calib_complete ,
    \asic/lsdram/msdram/io_dmi_cmd_ready ,
    \asic/lsdram/msdram/io_dmi_wr_data_rdy ,
    \asic/lsdram/msdram/io_dmi_rd_data_valid ,
    clock,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \asic/cpu/cpu/if_stage/fs_pc[31] ;
input \asic/cpu/cpu/if_stage/fs_pc[30] ;
input \asic/cpu/cpu/if_stage/fs_pc[29] ;
input \asic/cpu/cpu/if_stage/fs_pc[28] ;
input \asic/cpu/cpu/if_stage/fs_pc[27] ;
input \asic/cpu/cpu/if_stage/fs_pc[26] ;
input \asic/cpu/cpu/if_stage/fs_pc[25] ;
input \asic/cpu/cpu/if_stage/fs_pc[24] ;
input \asic/cpu/cpu/if_stage/fs_pc[23] ;
input \asic/cpu/cpu/if_stage/fs_pc[22] ;
input \asic/cpu/cpu/if_stage/fs_pc[21] ;
input \asic/cpu/cpu/if_stage/fs_pc[20] ;
input \asic/cpu/cpu/if_stage/fs_pc[19] ;
input \asic/cpu/cpu/if_stage/fs_pc[18] ;
input \asic/cpu/cpu/if_stage/fs_pc[17] ;
input \asic/cpu/cpu/if_stage/fs_pc[16] ;
input \asic/cpu/cpu/if_stage/fs_pc[15] ;
input \asic/cpu/cpu/if_stage/fs_pc[14] ;
input \asic/cpu/cpu/if_stage/fs_pc[13] ;
input \asic/cpu/cpu/if_stage/fs_pc[12] ;
input \asic/cpu/cpu/if_stage/fs_pc[11] ;
input \asic/cpu/cpu/if_stage/fs_pc[10] ;
input \asic/cpu/cpu/if_stage/fs_pc[9] ;
input \asic/cpu/cpu/if_stage/fs_pc[8] ;
input \asic/cpu/cpu/if_stage/fs_pc[7] ;
input \asic/cpu/cpu/if_stage/fs_pc[6] ;
input \asic/cpu/cpu/if_stage/fs_pc[5] ;
input \asic/cpu/cpu/if_stage/fs_pc[4] ;
input \asic/cpu/cpu/if_stage/fs_pc[3] ;
input \asic/cpu/cpu/if_stage/fs_pc[2] ;
input \asic/cpu/cpu/if_stage/fs_pc[1] ;
input \asic/cpu/cpu/if_stage/fs_pc[0] ;
input \asic/cpu/cpu/if_stage/fs_inst[31] ;
input \asic/cpu/cpu/if_stage/fs_inst[30] ;
input \asic/cpu/cpu/if_stage/fs_inst[29] ;
input \asic/cpu/cpu/if_stage/fs_inst[28] ;
input \asic/cpu/cpu/if_stage/fs_inst[27] ;
input \asic/cpu/cpu/if_stage/fs_inst[26] ;
input \asic/cpu/cpu/if_stage/fs_inst[25] ;
input \asic/cpu/cpu/if_stage/fs_inst[24] ;
input \asic/cpu/cpu/if_stage/fs_inst[23] ;
input \asic/cpu/cpu/if_stage/fs_inst[22] ;
input \asic/cpu/cpu/if_stage/fs_inst[21] ;
input \asic/cpu/cpu/if_stage/fs_inst[20] ;
input \asic/cpu/cpu/if_stage/fs_inst[19] ;
input \asic/cpu/cpu/if_stage/fs_inst[18] ;
input \asic/cpu/cpu/if_stage/fs_inst[17] ;
input \asic/cpu/cpu/if_stage/fs_inst[16] ;
input \asic/cpu/cpu/if_stage/fs_inst[15] ;
input \asic/cpu/cpu/if_stage/fs_inst[14] ;
input \asic/cpu/cpu/if_stage/fs_inst[13] ;
input \asic/cpu/cpu/if_stage/fs_inst[12] ;
input \asic/cpu/cpu/if_stage/fs_inst[11] ;
input \asic/cpu/cpu/if_stage/fs_inst[10] ;
input \asic/cpu/cpu/if_stage/fs_inst[9] ;
input \asic/cpu/cpu/if_stage/fs_inst[8] ;
input \asic/cpu/cpu/if_stage/fs_inst[7] ;
input \asic/cpu/cpu/if_stage/fs_inst[6] ;
input \asic/cpu/cpu/if_stage/fs_inst[5] ;
input \asic/cpu/cpu/if_stage/fs_inst[4] ;
input \asic/cpu/cpu/if_stage/fs_inst[3] ;
input \asic/cpu/cpu/if_stage/fs_inst[2] ;
input \asic/cpu/cpu/if_stage/fs_inst[1] ;
input \asic/cpu/cpu/if_stage/fs_inst[0] ;
input \asic/lsdram/msdram/io_in_awid[3] ;
input \asic/lsdram/msdram/io_in_awid[2] ;
input \asic/lsdram/msdram/io_in_awid[1] ;
input \asic/lsdram/msdram/io_in_awid[0] ;
input \asic/lsdram/msdram/io_in_awaddr[31] ;
input \asic/lsdram/msdram/io_in_awaddr[30] ;
input \asic/lsdram/msdram/io_in_awaddr[29] ;
input \asic/lsdram/msdram/io_in_awaddr[28] ;
input \asic/lsdram/msdram/io_in_awaddr[27] ;
input \asic/lsdram/msdram/io_in_awaddr[26] ;
input \asic/lsdram/msdram/io_in_awaddr[25] ;
input \asic/lsdram/msdram/io_in_awaddr[24] ;
input \asic/lsdram/msdram/io_in_awaddr[23] ;
input \asic/lsdram/msdram/io_in_awaddr[22] ;
input \asic/lsdram/msdram/io_in_awaddr[21] ;
input \asic/lsdram/msdram/io_in_awaddr[20] ;
input \asic/lsdram/msdram/io_in_awaddr[19] ;
input \asic/lsdram/msdram/io_in_awaddr[18] ;
input \asic/lsdram/msdram/io_in_awaddr[17] ;
input \asic/lsdram/msdram/io_in_awaddr[16] ;
input \asic/lsdram/msdram/io_in_awaddr[15] ;
input \asic/lsdram/msdram/io_in_awaddr[14] ;
input \asic/lsdram/msdram/io_in_awaddr[13] ;
input \asic/lsdram/msdram/io_in_awaddr[12] ;
input \asic/lsdram/msdram/io_in_awaddr[11] ;
input \asic/lsdram/msdram/io_in_awaddr[10] ;
input \asic/lsdram/msdram/io_in_awaddr[9] ;
input \asic/lsdram/msdram/io_in_awaddr[8] ;
input \asic/lsdram/msdram/io_in_awaddr[7] ;
input \asic/lsdram/msdram/io_in_awaddr[6] ;
input \asic/lsdram/msdram/io_in_awaddr[5] ;
input \asic/lsdram/msdram/io_in_awaddr[4] ;
input \asic/lsdram/msdram/io_in_awaddr[3] ;
input \asic/lsdram/msdram/io_in_awaddr[2] ;
input \asic/lsdram/msdram/io_in_awaddr[1] ;
input \asic/lsdram/msdram/io_in_awaddr[0] ;
input \asic/lsdram/msdram/io_in_awlen[7] ;
input \asic/lsdram/msdram/io_in_awlen[6] ;
input \asic/lsdram/msdram/io_in_awlen[5] ;
input \asic/lsdram/msdram/io_in_awlen[4] ;
input \asic/lsdram/msdram/io_in_awlen[3] ;
input \asic/lsdram/msdram/io_in_awlen[2] ;
input \asic/lsdram/msdram/io_in_awlen[1] ;
input \asic/lsdram/msdram/io_in_awlen[0] ;
input \asic/lsdram/msdram/io_in_awsize[2] ;
input \asic/lsdram/msdram/io_in_awsize[1] ;
input \asic/lsdram/msdram/io_in_awsize[0] ;
input \asic/lsdram/msdram/io_in_wdata[31] ;
input \asic/lsdram/msdram/io_in_wdata[30] ;
input \asic/lsdram/msdram/io_in_wdata[29] ;
input \asic/lsdram/msdram/io_in_wdata[28] ;
input \asic/lsdram/msdram/io_in_wdata[27] ;
input \asic/lsdram/msdram/io_in_wdata[26] ;
input \asic/lsdram/msdram/io_in_wdata[25] ;
input \asic/lsdram/msdram/io_in_wdata[24] ;
input \asic/lsdram/msdram/io_in_wdata[23] ;
input \asic/lsdram/msdram/io_in_wdata[22] ;
input \asic/lsdram/msdram/io_in_wdata[21] ;
input \asic/lsdram/msdram/io_in_wdata[20] ;
input \asic/lsdram/msdram/io_in_wdata[19] ;
input \asic/lsdram/msdram/io_in_wdata[18] ;
input \asic/lsdram/msdram/io_in_wdata[17] ;
input \asic/lsdram/msdram/io_in_wdata[16] ;
input \asic/lsdram/msdram/io_in_wdata[15] ;
input \asic/lsdram/msdram/io_in_wdata[14] ;
input \asic/lsdram/msdram/io_in_wdata[13] ;
input \asic/lsdram/msdram/io_in_wdata[12] ;
input \asic/lsdram/msdram/io_in_wdata[11] ;
input \asic/lsdram/msdram/io_in_wdata[10] ;
input \asic/lsdram/msdram/io_in_wdata[9] ;
input \asic/lsdram/msdram/io_in_wdata[8] ;
input \asic/lsdram/msdram/io_in_wdata[7] ;
input \asic/lsdram/msdram/io_in_wdata[6] ;
input \asic/lsdram/msdram/io_in_wdata[5] ;
input \asic/lsdram/msdram/io_in_wdata[4] ;
input \asic/lsdram/msdram/io_in_wdata[3] ;
input \asic/lsdram/msdram/io_in_wdata[2] ;
input \asic/lsdram/msdram/io_in_wdata[1] ;
input \asic/lsdram/msdram/io_in_wdata[0] ;
input \asic/lsdram/msdram/io_in_wstrb[3] ;
input \asic/lsdram/msdram/io_in_wstrb[2] ;
input \asic/lsdram/msdram/io_in_wstrb[1] ;
input \asic/lsdram/msdram/io_in_wstrb[0] ;
input \asic/lsdram/msdram/io_in_bid[3] ;
input \asic/lsdram/msdram/io_in_bid[2] ;
input \asic/lsdram/msdram/io_in_bid[1] ;
input \asic/lsdram/msdram/io_in_bid[0] ;
input \asic/lsdram/msdram/io_in_arid[3] ;
input \asic/lsdram/msdram/io_in_arid[2] ;
input \asic/lsdram/msdram/io_in_arid[1] ;
input \asic/lsdram/msdram/io_in_arid[0] ;
input \asic/lsdram/msdram/io_in_araddr[31] ;
input \asic/lsdram/msdram/io_in_araddr[30] ;
input \asic/lsdram/msdram/io_in_araddr[29] ;
input \asic/lsdram/msdram/io_in_araddr[28] ;
input \asic/lsdram/msdram/io_in_araddr[27] ;
input \asic/lsdram/msdram/io_in_araddr[26] ;
input \asic/lsdram/msdram/io_in_araddr[25] ;
input \asic/lsdram/msdram/io_in_araddr[24] ;
input \asic/lsdram/msdram/io_in_araddr[23] ;
input \asic/lsdram/msdram/io_in_araddr[22] ;
input \asic/lsdram/msdram/io_in_araddr[21] ;
input \asic/lsdram/msdram/io_in_araddr[20] ;
input \asic/lsdram/msdram/io_in_araddr[19] ;
input \asic/lsdram/msdram/io_in_araddr[18] ;
input \asic/lsdram/msdram/io_in_araddr[17] ;
input \asic/lsdram/msdram/io_in_araddr[16] ;
input \asic/lsdram/msdram/io_in_araddr[15] ;
input \asic/lsdram/msdram/io_in_araddr[14] ;
input \asic/lsdram/msdram/io_in_araddr[13] ;
input \asic/lsdram/msdram/io_in_araddr[12] ;
input \asic/lsdram/msdram/io_in_araddr[11] ;
input \asic/lsdram/msdram/io_in_araddr[10] ;
input \asic/lsdram/msdram/io_in_araddr[9] ;
input \asic/lsdram/msdram/io_in_araddr[8] ;
input \asic/lsdram/msdram/io_in_araddr[7] ;
input \asic/lsdram/msdram/io_in_araddr[6] ;
input \asic/lsdram/msdram/io_in_araddr[5] ;
input \asic/lsdram/msdram/io_in_araddr[4] ;
input \asic/lsdram/msdram/io_in_araddr[3] ;
input \asic/lsdram/msdram/io_in_araddr[2] ;
input \asic/lsdram/msdram/io_in_araddr[1] ;
input \asic/lsdram/msdram/io_in_araddr[0] ;
input \asic/lsdram/msdram/io_in_arlen[7] ;
input \asic/lsdram/msdram/io_in_arlen[6] ;
input \asic/lsdram/msdram/io_in_arlen[5] ;
input \asic/lsdram/msdram/io_in_arlen[4] ;
input \asic/lsdram/msdram/io_in_arlen[3] ;
input \asic/lsdram/msdram/io_in_arlen[2] ;
input \asic/lsdram/msdram/io_in_arlen[1] ;
input \asic/lsdram/msdram/io_in_arlen[0] ;
input \asic/lsdram/msdram/io_in_arsize[2] ;
input \asic/lsdram/msdram/io_in_arsize[1] ;
input \asic/lsdram/msdram/io_in_arsize[0] ;
input \asic/lsdram/msdram/io_in_rid[3] ;
input \asic/lsdram/msdram/io_in_rid[2] ;
input \asic/lsdram/msdram/io_in_rid[1] ;
input \asic/lsdram/msdram/io_in_rid[0] ;
input \asic/lsdram/msdram/io_in_rdata[31] ;
input \asic/lsdram/msdram/io_in_rdata[30] ;
input \asic/lsdram/msdram/io_in_rdata[29] ;
input \asic/lsdram/msdram/io_in_rdata[28] ;
input \asic/lsdram/msdram/io_in_rdata[27] ;
input \asic/lsdram/msdram/io_in_rdata[26] ;
input \asic/lsdram/msdram/io_in_rdata[25] ;
input \asic/lsdram/msdram/io_in_rdata[24] ;
input \asic/lsdram/msdram/io_in_rdata[23] ;
input \asic/lsdram/msdram/io_in_rdata[22] ;
input \asic/lsdram/msdram/io_in_rdata[21] ;
input \asic/lsdram/msdram/io_in_rdata[20] ;
input \asic/lsdram/msdram/io_in_rdata[19] ;
input \asic/lsdram/msdram/io_in_rdata[18] ;
input \asic/lsdram/msdram/io_in_rdata[17] ;
input \asic/lsdram/msdram/io_in_rdata[16] ;
input \asic/lsdram/msdram/io_in_rdata[15] ;
input \asic/lsdram/msdram/io_in_rdata[14] ;
input \asic/lsdram/msdram/io_in_rdata[13] ;
input \asic/lsdram/msdram/io_in_rdata[12] ;
input \asic/lsdram/msdram/io_in_rdata[11] ;
input \asic/lsdram/msdram/io_in_rdata[10] ;
input \asic/lsdram/msdram/io_in_rdata[9] ;
input \asic/lsdram/msdram/io_in_rdata[8] ;
input \asic/lsdram/msdram/io_in_rdata[7] ;
input \asic/lsdram/msdram/io_in_rdata[6] ;
input \asic/lsdram/msdram/io_in_rdata[5] ;
input \asic/lsdram/msdram/io_in_rdata[4] ;
input \asic/lsdram/msdram/io_in_rdata[3] ;
input \asic/lsdram/msdram/io_in_rdata[2] ;
input \asic/lsdram/msdram/io_in_rdata[1] ;
input \asic/lsdram/msdram/io_in_rdata[0] ;
input \asic/lsdram/msdram/io_dmi_cmd[2] ;
input \asic/lsdram/msdram/io_dmi_cmd[1] ;
input \asic/lsdram/msdram/io_dmi_cmd[0] ;
input \asic/lsdram/msdram/io_dmi_addr[28] ;
input \asic/lsdram/msdram/io_dmi_addr[27] ;
input \asic/lsdram/msdram/io_dmi_addr[26] ;
input \asic/lsdram/msdram/io_dmi_addr[25] ;
input \asic/lsdram/msdram/io_dmi_addr[24] ;
input \asic/lsdram/msdram/io_dmi_addr[23] ;
input \asic/lsdram/msdram/io_dmi_addr[22] ;
input \asic/lsdram/msdram/io_dmi_addr[21] ;
input \asic/lsdram/msdram/io_dmi_addr[20] ;
input \asic/lsdram/msdram/io_dmi_addr[19] ;
input \asic/lsdram/msdram/io_dmi_addr[18] ;
input \asic/lsdram/msdram/io_dmi_addr[17] ;
input \asic/lsdram/msdram/io_dmi_addr[16] ;
input \asic/lsdram/msdram/io_dmi_addr[15] ;
input \asic/lsdram/msdram/io_dmi_addr[14] ;
input \asic/lsdram/msdram/io_dmi_addr[13] ;
input \asic/lsdram/msdram/io_dmi_addr[12] ;
input \asic/lsdram/msdram/io_dmi_addr[11] ;
input \asic/lsdram/msdram/io_dmi_addr[10] ;
input \asic/lsdram/msdram/io_dmi_addr[9] ;
input \asic/lsdram/msdram/io_dmi_addr[8] ;
input \asic/lsdram/msdram/io_dmi_addr[7] ;
input \asic/lsdram/msdram/io_dmi_addr[6] ;
input \asic/lsdram/msdram/io_dmi_addr[5] ;
input \asic/lsdram/msdram/io_dmi_addr[4] ;
input \asic/lsdram/msdram/io_dmi_addr[3] ;
input \asic/lsdram/msdram/io_dmi_addr[2] ;
input \asic/lsdram/msdram/io_dmi_addr[1] ;
input \asic/lsdram/msdram/io_dmi_addr[0] ;
input \asic/lsdram/msdram/io_dmi_wr_data[255] ;
input \asic/lsdram/msdram/io_dmi_wr_data[254] ;
input \asic/lsdram/msdram/io_dmi_wr_data[253] ;
input \asic/lsdram/msdram/io_dmi_wr_data[252] ;
input \asic/lsdram/msdram/io_dmi_wr_data[251] ;
input \asic/lsdram/msdram/io_dmi_wr_data[250] ;
input \asic/lsdram/msdram/io_dmi_wr_data[249] ;
input \asic/lsdram/msdram/io_dmi_wr_data[248] ;
input \asic/lsdram/msdram/io_dmi_wr_data[247] ;
input \asic/lsdram/msdram/io_dmi_wr_data[246] ;
input \asic/lsdram/msdram/io_dmi_wr_data[245] ;
input \asic/lsdram/msdram/io_dmi_wr_data[244] ;
input \asic/lsdram/msdram/io_dmi_wr_data[243] ;
input \asic/lsdram/msdram/io_dmi_wr_data[242] ;
input \asic/lsdram/msdram/io_dmi_wr_data[241] ;
input \asic/lsdram/msdram/io_dmi_wr_data[240] ;
input \asic/lsdram/msdram/io_dmi_wr_data[239] ;
input \asic/lsdram/msdram/io_dmi_wr_data[238] ;
input \asic/lsdram/msdram/io_dmi_wr_data[237] ;
input \asic/lsdram/msdram/io_dmi_wr_data[236] ;
input \asic/lsdram/msdram/io_dmi_wr_data[235] ;
input \asic/lsdram/msdram/io_dmi_wr_data[234] ;
input \asic/lsdram/msdram/io_dmi_wr_data[233] ;
input \asic/lsdram/msdram/io_dmi_wr_data[232] ;
input \asic/lsdram/msdram/io_dmi_wr_data[231] ;
input \asic/lsdram/msdram/io_dmi_wr_data[230] ;
input \asic/lsdram/msdram/io_dmi_wr_data[229] ;
input \asic/lsdram/msdram/io_dmi_wr_data[228] ;
input \asic/lsdram/msdram/io_dmi_wr_data[227] ;
input \asic/lsdram/msdram/io_dmi_wr_data[226] ;
input \asic/lsdram/msdram/io_dmi_wr_data[225] ;
input \asic/lsdram/msdram/io_dmi_wr_data[224] ;
input \asic/lsdram/msdram/io_dmi_wr_data[223] ;
input \asic/lsdram/msdram/io_dmi_wr_data[222] ;
input \asic/lsdram/msdram/io_dmi_wr_data[221] ;
input \asic/lsdram/msdram/io_dmi_wr_data[220] ;
input \asic/lsdram/msdram/io_dmi_wr_data[219] ;
input \asic/lsdram/msdram/io_dmi_wr_data[218] ;
input \asic/lsdram/msdram/io_dmi_wr_data[217] ;
input \asic/lsdram/msdram/io_dmi_wr_data[216] ;
input \asic/lsdram/msdram/io_dmi_wr_data[215] ;
input \asic/lsdram/msdram/io_dmi_wr_data[214] ;
input \asic/lsdram/msdram/io_dmi_wr_data[213] ;
input \asic/lsdram/msdram/io_dmi_wr_data[212] ;
input \asic/lsdram/msdram/io_dmi_wr_data[211] ;
input \asic/lsdram/msdram/io_dmi_wr_data[210] ;
input \asic/lsdram/msdram/io_dmi_wr_data[209] ;
input \asic/lsdram/msdram/io_dmi_wr_data[208] ;
input \asic/lsdram/msdram/io_dmi_wr_data[207] ;
input \asic/lsdram/msdram/io_dmi_wr_data[206] ;
input \asic/lsdram/msdram/io_dmi_wr_data[205] ;
input \asic/lsdram/msdram/io_dmi_wr_data[204] ;
input \asic/lsdram/msdram/io_dmi_wr_data[203] ;
input \asic/lsdram/msdram/io_dmi_wr_data[202] ;
input \asic/lsdram/msdram/io_dmi_wr_data[201] ;
input \asic/lsdram/msdram/io_dmi_wr_data[200] ;
input \asic/lsdram/msdram/io_dmi_wr_data[199] ;
input \asic/lsdram/msdram/io_dmi_wr_data[198] ;
input \asic/lsdram/msdram/io_dmi_wr_data[197] ;
input \asic/lsdram/msdram/io_dmi_wr_data[196] ;
input \asic/lsdram/msdram/io_dmi_wr_data[195] ;
input \asic/lsdram/msdram/io_dmi_wr_data[194] ;
input \asic/lsdram/msdram/io_dmi_wr_data[193] ;
input \asic/lsdram/msdram/io_dmi_wr_data[192] ;
input \asic/lsdram/msdram/io_dmi_wr_data[191] ;
input \asic/lsdram/msdram/io_dmi_wr_data[190] ;
input \asic/lsdram/msdram/io_dmi_wr_data[189] ;
input \asic/lsdram/msdram/io_dmi_wr_data[188] ;
input \asic/lsdram/msdram/io_dmi_wr_data[187] ;
input \asic/lsdram/msdram/io_dmi_wr_data[186] ;
input \asic/lsdram/msdram/io_dmi_wr_data[185] ;
input \asic/lsdram/msdram/io_dmi_wr_data[184] ;
input \asic/lsdram/msdram/io_dmi_wr_data[183] ;
input \asic/lsdram/msdram/io_dmi_wr_data[182] ;
input \asic/lsdram/msdram/io_dmi_wr_data[181] ;
input \asic/lsdram/msdram/io_dmi_wr_data[180] ;
input \asic/lsdram/msdram/io_dmi_wr_data[179] ;
input \asic/lsdram/msdram/io_dmi_wr_data[178] ;
input \asic/lsdram/msdram/io_dmi_wr_data[177] ;
input \asic/lsdram/msdram/io_dmi_wr_data[176] ;
input \asic/lsdram/msdram/io_dmi_wr_data[175] ;
input \asic/lsdram/msdram/io_dmi_wr_data[174] ;
input \asic/lsdram/msdram/io_dmi_wr_data[173] ;
input \asic/lsdram/msdram/io_dmi_wr_data[172] ;
input \asic/lsdram/msdram/io_dmi_wr_data[171] ;
input \asic/lsdram/msdram/io_dmi_wr_data[170] ;
input \asic/lsdram/msdram/io_dmi_wr_data[169] ;
input \asic/lsdram/msdram/io_dmi_wr_data[168] ;
input \asic/lsdram/msdram/io_dmi_wr_data[167] ;
input \asic/lsdram/msdram/io_dmi_wr_data[166] ;
input \asic/lsdram/msdram/io_dmi_wr_data[165] ;
input \asic/lsdram/msdram/io_dmi_wr_data[164] ;
input \asic/lsdram/msdram/io_dmi_wr_data[163] ;
input \asic/lsdram/msdram/io_dmi_wr_data[162] ;
input \asic/lsdram/msdram/io_dmi_wr_data[161] ;
input \asic/lsdram/msdram/io_dmi_wr_data[160] ;
input \asic/lsdram/msdram/io_dmi_wr_data[159] ;
input \asic/lsdram/msdram/io_dmi_wr_data[158] ;
input \asic/lsdram/msdram/io_dmi_wr_data[157] ;
input \asic/lsdram/msdram/io_dmi_wr_data[156] ;
input \asic/lsdram/msdram/io_dmi_wr_data[155] ;
input \asic/lsdram/msdram/io_dmi_wr_data[154] ;
input \asic/lsdram/msdram/io_dmi_wr_data[153] ;
input \asic/lsdram/msdram/io_dmi_wr_data[152] ;
input \asic/lsdram/msdram/io_dmi_wr_data[151] ;
input \asic/lsdram/msdram/io_dmi_wr_data[150] ;
input \asic/lsdram/msdram/io_dmi_wr_data[149] ;
input \asic/lsdram/msdram/io_dmi_wr_data[148] ;
input \asic/lsdram/msdram/io_dmi_wr_data[147] ;
input \asic/lsdram/msdram/io_dmi_wr_data[146] ;
input \asic/lsdram/msdram/io_dmi_wr_data[145] ;
input \asic/lsdram/msdram/io_dmi_wr_data[144] ;
input \asic/lsdram/msdram/io_dmi_wr_data[143] ;
input \asic/lsdram/msdram/io_dmi_wr_data[142] ;
input \asic/lsdram/msdram/io_dmi_wr_data[141] ;
input \asic/lsdram/msdram/io_dmi_wr_data[140] ;
input \asic/lsdram/msdram/io_dmi_wr_data[139] ;
input \asic/lsdram/msdram/io_dmi_wr_data[138] ;
input \asic/lsdram/msdram/io_dmi_wr_data[137] ;
input \asic/lsdram/msdram/io_dmi_wr_data[136] ;
input \asic/lsdram/msdram/io_dmi_wr_data[135] ;
input \asic/lsdram/msdram/io_dmi_wr_data[134] ;
input \asic/lsdram/msdram/io_dmi_wr_data[133] ;
input \asic/lsdram/msdram/io_dmi_wr_data[132] ;
input \asic/lsdram/msdram/io_dmi_wr_data[131] ;
input \asic/lsdram/msdram/io_dmi_wr_data[130] ;
input \asic/lsdram/msdram/io_dmi_wr_data[129] ;
input \asic/lsdram/msdram/io_dmi_wr_data[128] ;
input \asic/lsdram/msdram/io_dmi_wr_data[127] ;
input \asic/lsdram/msdram/io_dmi_wr_data[126] ;
input \asic/lsdram/msdram/io_dmi_wr_data[125] ;
input \asic/lsdram/msdram/io_dmi_wr_data[124] ;
input \asic/lsdram/msdram/io_dmi_wr_data[123] ;
input \asic/lsdram/msdram/io_dmi_wr_data[122] ;
input \asic/lsdram/msdram/io_dmi_wr_data[121] ;
input \asic/lsdram/msdram/io_dmi_wr_data[120] ;
input \asic/lsdram/msdram/io_dmi_wr_data[119] ;
input \asic/lsdram/msdram/io_dmi_wr_data[118] ;
input \asic/lsdram/msdram/io_dmi_wr_data[117] ;
input \asic/lsdram/msdram/io_dmi_wr_data[116] ;
input \asic/lsdram/msdram/io_dmi_wr_data[115] ;
input \asic/lsdram/msdram/io_dmi_wr_data[114] ;
input \asic/lsdram/msdram/io_dmi_wr_data[113] ;
input \asic/lsdram/msdram/io_dmi_wr_data[112] ;
input \asic/lsdram/msdram/io_dmi_wr_data[111] ;
input \asic/lsdram/msdram/io_dmi_wr_data[110] ;
input \asic/lsdram/msdram/io_dmi_wr_data[109] ;
input \asic/lsdram/msdram/io_dmi_wr_data[108] ;
input \asic/lsdram/msdram/io_dmi_wr_data[107] ;
input \asic/lsdram/msdram/io_dmi_wr_data[106] ;
input \asic/lsdram/msdram/io_dmi_wr_data[105] ;
input \asic/lsdram/msdram/io_dmi_wr_data[104] ;
input \asic/lsdram/msdram/io_dmi_wr_data[103] ;
input \asic/lsdram/msdram/io_dmi_wr_data[102] ;
input \asic/lsdram/msdram/io_dmi_wr_data[101] ;
input \asic/lsdram/msdram/io_dmi_wr_data[100] ;
input \asic/lsdram/msdram/io_dmi_wr_data[99] ;
input \asic/lsdram/msdram/io_dmi_wr_data[98] ;
input \asic/lsdram/msdram/io_dmi_wr_data[97] ;
input \asic/lsdram/msdram/io_dmi_wr_data[96] ;
input \asic/lsdram/msdram/io_dmi_wr_data[95] ;
input \asic/lsdram/msdram/io_dmi_wr_data[94] ;
input \asic/lsdram/msdram/io_dmi_wr_data[93] ;
input \asic/lsdram/msdram/io_dmi_wr_data[92] ;
input \asic/lsdram/msdram/io_dmi_wr_data[91] ;
input \asic/lsdram/msdram/io_dmi_wr_data[90] ;
input \asic/lsdram/msdram/io_dmi_wr_data[89] ;
input \asic/lsdram/msdram/io_dmi_wr_data[88] ;
input \asic/lsdram/msdram/io_dmi_wr_data[87] ;
input \asic/lsdram/msdram/io_dmi_wr_data[86] ;
input \asic/lsdram/msdram/io_dmi_wr_data[85] ;
input \asic/lsdram/msdram/io_dmi_wr_data[84] ;
input \asic/lsdram/msdram/io_dmi_wr_data[83] ;
input \asic/lsdram/msdram/io_dmi_wr_data[82] ;
input \asic/lsdram/msdram/io_dmi_wr_data[81] ;
input \asic/lsdram/msdram/io_dmi_wr_data[80] ;
input \asic/lsdram/msdram/io_dmi_wr_data[79] ;
input \asic/lsdram/msdram/io_dmi_wr_data[78] ;
input \asic/lsdram/msdram/io_dmi_wr_data[77] ;
input \asic/lsdram/msdram/io_dmi_wr_data[76] ;
input \asic/lsdram/msdram/io_dmi_wr_data[75] ;
input \asic/lsdram/msdram/io_dmi_wr_data[74] ;
input \asic/lsdram/msdram/io_dmi_wr_data[73] ;
input \asic/lsdram/msdram/io_dmi_wr_data[72] ;
input \asic/lsdram/msdram/io_dmi_wr_data[71] ;
input \asic/lsdram/msdram/io_dmi_wr_data[70] ;
input \asic/lsdram/msdram/io_dmi_wr_data[69] ;
input \asic/lsdram/msdram/io_dmi_wr_data[68] ;
input \asic/lsdram/msdram/io_dmi_wr_data[67] ;
input \asic/lsdram/msdram/io_dmi_wr_data[66] ;
input \asic/lsdram/msdram/io_dmi_wr_data[65] ;
input \asic/lsdram/msdram/io_dmi_wr_data[64] ;
input \asic/lsdram/msdram/io_dmi_wr_data[63] ;
input \asic/lsdram/msdram/io_dmi_wr_data[62] ;
input \asic/lsdram/msdram/io_dmi_wr_data[61] ;
input \asic/lsdram/msdram/io_dmi_wr_data[60] ;
input \asic/lsdram/msdram/io_dmi_wr_data[59] ;
input \asic/lsdram/msdram/io_dmi_wr_data[58] ;
input \asic/lsdram/msdram/io_dmi_wr_data[57] ;
input \asic/lsdram/msdram/io_dmi_wr_data[56] ;
input \asic/lsdram/msdram/io_dmi_wr_data[55] ;
input \asic/lsdram/msdram/io_dmi_wr_data[54] ;
input \asic/lsdram/msdram/io_dmi_wr_data[53] ;
input \asic/lsdram/msdram/io_dmi_wr_data[52] ;
input \asic/lsdram/msdram/io_dmi_wr_data[51] ;
input \asic/lsdram/msdram/io_dmi_wr_data[50] ;
input \asic/lsdram/msdram/io_dmi_wr_data[49] ;
input \asic/lsdram/msdram/io_dmi_wr_data[48] ;
input \asic/lsdram/msdram/io_dmi_wr_data[47] ;
input \asic/lsdram/msdram/io_dmi_wr_data[46] ;
input \asic/lsdram/msdram/io_dmi_wr_data[45] ;
input \asic/lsdram/msdram/io_dmi_wr_data[44] ;
input \asic/lsdram/msdram/io_dmi_wr_data[43] ;
input \asic/lsdram/msdram/io_dmi_wr_data[42] ;
input \asic/lsdram/msdram/io_dmi_wr_data[41] ;
input \asic/lsdram/msdram/io_dmi_wr_data[40] ;
input \asic/lsdram/msdram/io_dmi_wr_data[39] ;
input \asic/lsdram/msdram/io_dmi_wr_data[38] ;
input \asic/lsdram/msdram/io_dmi_wr_data[37] ;
input \asic/lsdram/msdram/io_dmi_wr_data[36] ;
input \asic/lsdram/msdram/io_dmi_wr_data[35] ;
input \asic/lsdram/msdram/io_dmi_wr_data[34] ;
input \asic/lsdram/msdram/io_dmi_wr_data[33] ;
input \asic/lsdram/msdram/io_dmi_wr_data[32] ;
input \asic/lsdram/msdram/io_dmi_wr_data[31] ;
input \asic/lsdram/msdram/io_dmi_wr_data[30] ;
input \asic/lsdram/msdram/io_dmi_wr_data[29] ;
input \asic/lsdram/msdram/io_dmi_wr_data[28] ;
input \asic/lsdram/msdram/io_dmi_wr_data[27] ;
input \asic/lsdram/msdram/io_dmi_wr_data[26] ;
input \asic/lsdram/msdram/io_dmi_wr_data[25] ;
input \asic/lsdram/msdram/io_dmi_wr_data[24] ;
input \asic/lsdram/msdram/io_dmi_wr_data[23] ;
input \asic/lsdram/msdram/io_dmi_wr_data[22] ;
input \asic/lsdram/msdram/io_dmi_wr_data[21] ;
input \asic/lsdram/msdram/io_dmi_wr_data[20] ;
input \asic/lsdram/msdram/io_dmi_wr_data[19] ;
input \asic/lsdram/msdram/io_dmi_wr_data[18] ;
input \asic/lsdram/msdram/io_dmi_wr_data[17] ;
input \asic/lsdram/msdram/io_dmi_wr_data[16] ;
input \asic/lsdram/msdram/io_dmi_wr_data[15] ;
input \asic/lsdram/msdram/io_dmi_wr_data[14] ;
input \asic/lsdram/msdram/io_dmi_wr_data[13] ;
input \asic/lsdram/msdram/io_dmi_wr_data[12] ;
input \asic/lsdram/msdram/io_dmi_wr_data[11] ;
input \asic/lsdram/msdram/io_dmi_wr_data[10] ;
input \asic/lsdram/msdram/io_dmi_wr_data[9] ;
input \asic/lsdram/msdram/io_dmi_wr_data[8] ;
input \asic/lsdram/msdram/io_dmi_wr_data[7] ;
input \asic/lsdram/msdram/io_dmi_wr_data[6] ;
input \asic/lsdram/msdram/io_dmi_wr_data[5] ;
input \asic/lsdram/msdram/io_dmi_wr_data[4] ;
input \asic/lsdram/msdram/io_dmi_wr_data[3] ;
input \asic/lsdram/msdram/io_dmi_wr_data[2] ;
input \asic/lsdram/msdram/io_dmi_wr_data[1] ;
input \asic/lsdram/msdram/io_dmi_wr_data[0] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[31] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[30] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[29] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[28] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[27] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[26] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[25] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[24] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[23] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[22] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[21] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[20] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[19] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[18] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[17] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[16] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[15] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[14] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[13] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[12] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[11] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[10] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[9] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[8] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[7] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[6] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[5] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[4] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[3] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[2] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[1] ;
input \asic/lsdram/msdram/io_dmi_wr_data_mask[0] ;
input \asic/lsdram/msdram/io_dmi_rd_data[255] ;
input \asic/lsdram/msdram/io_dmi_rd_data[254] ;
input \asic/lsdram/msdram/io_dmi_rd_data[253] ;
input \asic/lsdram/msdram/io_dmi_rd_data[252] ;
input \asic/lsdram/msdram/io_dmi_rd_data[251] ;
input \asic/lsdram/msdram/io_dmi_rd_data[250] ;
input \asic/lsdram/msdram/io_dmi_rd_data[249] ;
input \asic/lsdram/msdram/io_dmi_rd_data[248] ;
input \asic/lsdram/msdram/io_dmi_rd_data[247] ;
input \asic/lsdram/msdram/io_dmi_rd_data[246] ;
input \asic/lsdram/msdram/io_dmi_rd_data[245] ;
input \asic/lsdram/msdram/io_dmi_rd_data[244] ;
input \asic/lsdram/msdram/io_dmi_rd_data[243] ;
input \asic/lsdram/msdram/io_dmi_rd_data[242] ;
input \asic/lsdram/msdram/io_dmi_rd_data[241] ;
input \asic/lsdram/msdram/io_dmi_rd_data[240] ;
input \asic/lsdram/msdram/io_dmi_rd_data[239] ;
input \asic/lsdram/msdram/io_dmi_rd_data[238] ;
input \asic/lsdram/msdram/io_dmi_rd_data[237] ;
input \asic/lsdram/msdram/io_dmi_rd_data[236] ;
input \asic/lsdram/msdram/io_dmi_rd_data[235] ;
input \asic/lsdram/msdram/io_dmi_rd_data[234] ;
input \asic/lsdram/msdram/io_dmi_rd_data[233] ;
input \asic/lsdram/msdram/io_dmi_rd_data[232] ;
input \asic/lsdram/msdram/io_dmi_rd_data[231] ;
input \asic/lsdram/msdram/io_dmi_rd_data[230] ;
input \asic/lsdram/msdram/io_dmi_rd_data[229] ;
input \asic/lsdram/msdram/io_dmi_rd_data[228] ;
input \asic/lsdram/msdram/io_dmi_rd_data[227] ;
input \asic/lsdram/msdram/io_dmi_rd_data[226] ;
input \asic/lsdram/msdram/io_dmi_rd_data[225] ;
input \asic/lsdram/msdram/io_dmi_rd_data[224] ;
input \asic/lsdram/msdram/io_dmi_rd_data[223] ;
input \asic/lsdram/msdram/io_dmi_rd_data[222] ;
input \asic/lsdram/msdram/io_dmi_rd_data[221] ;
input \asic/lsdram/msdram/io_dmi_rd_data[220] ;
input \asic/lsdram/msdram/io_dmi_rd_data[219] ;
input \asic/lsdram/msdram/io_dmi_rd_data[218] ;
input \asic/lsdram/msdram/io_dmi_rd_data[217] ;
input \asic/lsdram/msdram/io_dmi_rd_data[216] ;
input \asic/lsdram/msdram/io_dmi_rd_data[215] ;
input \asic/lsdram/msdram/io_dmi_rd_data[214] ;
input \asic/lsdram/msdram/io_dmi_rd_data[213] ;
input \asic/lsdram/msdram/io_dmi_rd_data[212] ;
input \asic/lsdram/msdram/io_dmi_rd_data[211] ;
input \asic/lsdram/msdram/io_dmi_rd_data[210] ;
input \asic/lsdram/msdram/io_dmi_rd_data[209] ;
input \asic/lsdram/msdram/io_dmi_rd_data[208] ;
input \asic/lsdram/msdram/io_dmi_rd_data[207] ;
input \asic/lsdram/msdram/io_dmi_rd_data[206] ;
input \asic/lsdram/msdram/io_dmi_rd_data[205] ;
input \asic/lsdram/msdram/io_dmi_rd_data[204] ;
input \asic/lsdram/msdram/io_dmi_rd_data[203] ;
input \asic/lsdram/msdram/io_dmi_rd_data[202] ;
input \asic/lsdram/msdram/io_dmi_rd_data[201] ;
input \asic/lsdram/msdram/io_dmi_rd_data[200] ;
input \asic/lsdram/msdram/io_dmi_rd_data[199] ;
input \asic/lsdram/msdram/io_dmi_rd_data[198] ;
input \asic/lsdram/msdram/io_dmi_rd_data[197] ;
input \asic/lsdram/msdram/io_dmi_rd_data[196] ;
input \asic/lsdram/msdram/io_dmi_rd_data[195] ;
input \asic/lsdram/msdram/io_dmi_rd_data[194] ;
input \asic/lsdram/msdram/io_dmi_rd_data[193] ;
input \asic/lsdram/msdram/io_dmi_rd_data[192] ;
input \asic/lsdram/msdram/io_dmi_rd_data[191] ;
input \asic/lsdram/msdram/io_dmi_rd_data[190] ;
input \asic/lsdram/msdram/io_dmi_rd_data[189] ;
input \asic/lsdram/msdram/io_dmi_rd_data[188] ;
input \asic/lsdram/msdram/io_dmi_rd_data[187] ;
input \asic/lsdram/msdram/io_dmi_rd_data[186] ;
input \asic/lsdram/msdram/io_dmi_rd_data[185] ;
input \asic/lsdram/msdram/io_dmi_rd_data[184] ;
input \asic/lsdram/msdram/io_dmi_rd_data[183] ;
input \asic/lsdram/msdram/io_dmi_rd_data[182] ;
input \asic/lsdram/msdram/io_dmi_rd_data[181] ;
input \asic/lsdram/msdram/io_dmi_rd_data[180] ;
input \asic/lsdram/msdram/io_dmi_rd_data[179] ;
input \asic/lsdram/msdram/io_dmi_rd_data[178] ;
input \asic/lsdram/msdram/io_dmi_rd_data[177] ;
input \asic/lsdram/msdram/io_dmi_rd_data[176] ;
input \asic/lsdram/msdram/io_dmi_rd_data[175] ;
input \asic/lsdram/msdram/io_dmi_rd_data[174] ;
input \asic/lsdram/msdram/io_dmi_rd_data[173] ;
input \asic/lsdram/msdram/io_dmi_rd_data[172] ;
input \asic/lsdram/msdram/io_dmi_rd_data[171] ;
input \asic/lsdram/msdram/io_dmi_rd_data[170] ;
input \asic/lsdram/msdram/io_dmi_rd_data[169] ;
input \asic/lsdram/msdram/io_dmi_rd_data[168] ;
input \asic/lsdram/msdram/io_dmi_rd_data[167] ;
input \asic/lsdram/msdram/io_dmi_rd_data[166] ;
input \asic/lsdram/msdram/io_dmi_rd_data[165] ;
input \asic/lsdram/msdram/io_dmi_rd_data[164] ;
input \asic/lsdram/msdram/io_dmi_rd_data[163] ;
input \asic/lsdram/msdram/io_dmi_rd_data[162] ;
input \asic/lsdram/msdram/io_dmi_rd_data[161] ;
input \asic/lsdram/msdram/io_dmi_rd_data[160] ;
input \asic/lsdram/msdram/io_dmi_rd_data[159] ;
input \asic/lsdram/msdram/io_dmi_rd_data[158] ;
input \asic/lsdram/msdram/io_dmi_rd_data[157] ;
input \asic/lsdram/msdram/io_dmi_rd_data[156] ;
input \asic/lsdram/msdram/io_dmi_rd_data[155] ;
input \asic/lsdram/msdram/io_dmi_rd_data[154] ;
input \asic/lsdram/msdram/io_dmi_rd_data[153] ;
input \asic/lsdram/msdram/io_dmi_rd_data[152] ;
input \asic/lsdram/msdram/io_dmi_rd_data[151] ;
input \asic/lsdram/msdram/io_dmi_rd_data[150] ;
input \asic/lsdram/msdram/io_dmi_rd_data[149] ;
input \asic/lsdram/msdram/io_dmi_rd_data[148] ;
input \asic/lsdram/msdram/io_dmi_rd_data[147] ;
input \asic/lsdram/msdram/io_dmi_rd_data[146] ;
input \asic/lsdram/msdram/io_dmi_rd_data[145] ;
input \asic/lsdram/msdram/io_dmi_rd_data[144] ;
input \asic/lsdram/msdram/io_dmi_rd_data[143] ;
input \asic/lsdram/msdram/io_dmi_rd_data[142] ;
input \asic/lsdram/msdram/io_dmi_rd_data[141] ;
input \asic/lsdram/msdram/io_dmi_rd_data[140] ;
input \asic/lsdram/msdram/io_dmi_rd_data[139] ;
input \asic/lsdram/msdram/io_dmi_rd_data[138] ;
input \asic/lsdram/msdram/io_dmi_rd_data[137] ;
input \asic/lsdram/msdram/io_dmi_rd_data[136] ;
input \asic/lsdram/msdram/io_dmi_rd_data[135] ;
input \asic/lsdram/msdram/io_dmi_rd_data[134] ;
input \asic/lsdram/msdram/io_dmi_rd_data[133] ;
input \asic/lsdram/msdram/io_dmi_rd_data[132] ;
input \asic/lsdram/msdram/io_dmi_rd_data[131] ;
input \asic/lsdram/msdram/io_dmi_rd_data[130] ;
input \asic/lsdram/msdram/io_dmi_rd_data[129] ;
input \asic/lsdram/msdram/io_dmi_rd_data[128] ;
input \asic/lsdram/msdram/io_dmi_rd_data[127] ;
input \asic/lsdram/msdram/io_dmi_rd_data[126] ;
input \asic/lsdram/msdram/io_dmi_rd_data[125] ;
input \asic/lsdram/msdram/io_dmi_rd_data[124] ;
input \asic/lsdram/msdram/io_dmi_rd_data[123] ;
input \asic/lsdram/msdram/io_dmi_rd_data[122] ;
input \asic/lsdram/msdram/io_dmi_rd_data[121] ;
input \asic/lsdram/msdram/io_dmi_rd_data[120] ;
input \asic/lsdram/msdram/io_dmi_rd_data[119] ;
input \asic/lsdram/msdram/io_dmi_rd_data[118] ;
input \asic/lsdram/msdram/io_dmi_rd_data[117] ;
input \asic/lsdram/msdram/io_dmi_rd_data[116] ;
input \asic/lsdram/msdram/io_dmi_rd_data[115] ;
input \asic/lsdram/msdram/io_dmi_rd_data[114] ;
input \asic/lsdram/msdram/io_dmi_rd_data[113] ;
input \asic/lsdram/msdram/io_dmi_rd_data[112] ;
input \asic/lsdram/msdram/io_dmi_rd_data[111] ;
input \asic/lsdram/msdram/io_dmi_rd_data[110] ;
input \asic/lsdram/msdram/io_dmi_rd_data[109] ;
input \asic/lsdram/msdram/io_dmi_rd_data[108] ;
input \asic/lsdram/msdram/io_dmi_rd_data[107] ;
input \asic/lsdram/msdram/io_dmi_rd_data[106] ;
input \asic/lsdram/msdram/io_dmi_rd_data[105] ;
input \asic/lsdram/msdram/io_dmi_rd_data[104] ;
input \asic/lsdram/msdram/io_dmi_rd_data[103] ;
input \asic/lsdram/msdram/io_dmi_rd_data[102] ;
input \asic/lsdram/msdram/io_dmi_rd_data[101] ;
input \asic/lsdram/msdram/io_dmi_rd_data[100] ;
input \asic/lsdram/msdram/io_dmi_rd_data[99] ;
input \asic/lsdram/msdram/io_dmi_rd_data[98] ;
input \asic/lsdram/msdram/io_dmi_rd_data[97] ;
input \asic/lsdram/msdram/io_dmi_rd_data[96] ;
input \asic/lsdram/msdram/io_dmi_rd_data[95] ;
input \asic/lsdram/msdram/io_dmi_rd_data[94] ;
input \asic/lsdram/msdram/io_dmi_rd_data[93] ;
input \asic/lsdram/msdram/io_dmi_rd_data[92] ;
input \asic/lsdram/msdram/io_dmi_rd_data[91] ;
input \asic/lsdram/msdram/io_dmi_rd_data[90] ;
input \asic/lsdram/msdram/io_dmi_rd_data[89] ;
input \asic/lsdram/msdram/io_dmi_rd_data[88] ;
input \asic/lsdram/msdram/io_dmi_rd_data[87] ;
input \asic/lsdram/msdram/io_dmi_rd_data[86] ;
input \asic/lsdram/msdram/io_dmi_rd_data[85] ;
input \asic/lsdram/msdram/io_dmi_rd_data[84] ;
input \asic/lsdram/msdram/io_dmi_rd_data[83] ;
input \asic/lsdram/msdram/io_dmi_rd_data[82] ;
input \asic/lsdram/msdram/io_dmi_rd_data[81] ;
input \asic/lsdram/msdram/io_dmi_rd_data[80] ;
input \asic/lsdram/msdram/io_dmi_rd_data[79] ;
input \asic/lsdram/msdram/io_dmi_rd_data[78] ;
input \asic/lsdram/msdram/io_dmi_rd_data[77] ;
input \asic/lsdram/msdram/io_dmi_rd_data[76] ;
input \asic/lsdram/msdram/io_dmi_rd_data[75] ;
input \asic/lsdram/msdram/io_dmi_rd_data[74] ;
input \asic/lsdram/msdram/io_dmi_rd_data[73] ;
input \asic/lsdram/msdram/io_dmi_rd_data[72] ;
input \asic/lsdram/msdram/io_dmi_rd_data[71] ;
input \asic/lsdram/msdram/io_dmi_rd_data[70] ;
input \asic/lsdram/msdram/io_dmi_rd_data[69] ;
input \asic/lsdram/msdram/io_dmi_rd_data[68] ;
input \asic/lsdram/msdram/io_dmi_rd_data[67] ;
input \asic/lsdram/msdram/io_dmi_rd_data[66] ;
input \asic/lsdram/msdram/io_dmi_rd_data[65] ;
input \asic/lsdram/msdram/io_dmi_rd_data[64] ;
input \asic/lsdram/msdram/io_dmi_rd_data[63] ;
input \asic/lsdram/msdram/io_dmi_rd_data[62] ;
input \asic/lsdram/msdram/io_dmi_rd_data[61] ;
input \asic/lsdram/msdram/io_dmi_rd_data[60] ;
input \asic/lsdram/msdram/io_dmi_rd_data[59] ;
input \asic/lsdram/msdram/io_dmi_rd_data[58] ;
input \asic/lsdram/msdram/io_dmi_rd_data[57] ;
input \asic/lsdram/msdram/io_dmi_rd_data[56] ;
input \asic/lsdram/msdram/io_dmi_rd_data[55] ;
input \asic/lsdram/msdram/io_dmi_rd_data[54] ;
input \asic/lsdram/msdram/io_dmi_rd_data[53] ;
input \asic/lsdram/msdram/io_dmi_rd_data[52] ;
input \asic/lsdram/msdram/io_dmi_rd_data[51] ;
input \asic/lsdram/msdram/io_dmi_rd_data[50] ;
input \asic/lsdram/msdram/io_dmi_rd_data[49] ;
input \asic/lsdram/msdram/io_dmi_rd_data[48] ;
input \asic/lsdram/msdram/io_dmi_rd_data[47] ;
input \asic/lsdram/msdram/io_dmi_rd_data[46] ;
input \asic/lsdram/msdram/io_dmi_rd_data[45] ;
input \asic/lsdram/msdram/io_dmi_rd_data[44] ;
input \asic/lsdram/msdram/io_dmi_rd_data[43] ;
input \asic/lsdram/msdram/io_dmi_rd_data[42] ;
input \asic/lsdram/msdram/io_dmi_rd_data[41] ;
input \asic/lsdram/msdram/io_dmi_rd_data[40] ;
input \asic/lsdram/msdram/io_dmi_rd_data[39] ;
input \asic/lsdram/msdram/io_dmi_rd_data[38] ;
input \asic/lsdram/msdram/io_dmi_rd_data[37] ;
input \asic/lsdram/msdram/io_dmi_rd_data[36] ;
input \asic/lsdram/msdram/io_dmi_rd_data[35] ;
input \asic/lsdram/msdram/io_dmi_rd_data[34] ;
input \asic/lsdram/msdram/io_dmi_rd_data[33] ;
input \asic/lsdram/msdram/io_dmi_rd_data[32] ;
input \asic/lsdram/msdram/io_dmi_rd_data[31] ;
input \asic/lsdram/msdram/io_dmi_rd_data[30] ;
input \asic/lsdram/msdram/io_dmi_rd_data[29] ;
input \asic/lsdram/msdram/io_dmi_rd_data[28] ;
input \asic/lsdram/msdram/io_dmi_rd_data[27] ;
input \asic/lsdram/msdram/io_dmi_rd_data[26] ;
input \asic/lsdram/msdram/io_dmi_rd_data[25] ;
input \asic/lsdram/msdram/io_dmi_rd_data[24] ;
input \asic/lsdram/msdram/io_dmi_rd_data[23] ;
input \asic/lsdram/msdram/io_dmi_rd_data[22] ;
input \asic/lsdram/msdram/io_dmi_rd_data[21] ;
input \asic/lsdram/msdram/io_dmi_rd_data[20] ;
input \asic/lsdram/msdram/io_dmi_rd_data[19] ;
input \asic/lsdram/msdram/io_dmi_rd_data[18] ;
input \asic/lsdram/msdram/io_dmi_rd_data[17] ;
input \asic/lsdram/msdram/io_dmi_rd_data[16] ;
input \asic/lsdram/msdram/io_dmi_rd_data[15] ;
input \asic/lsdram/msdram/io_dmi_rd_data[14] ;
input \asic/lsdram/msdram/io_dmi_rd_data[13] ;
input \asic/lsdram/msdram/io_dmi_rd_data[12] ;
input \asic/lsdram/msdram/io_dmi_rd_data[11] ;
input \asic/lsdram/msdram/io_dmi_rd_data[10] ;
input \asic/lsdram/msdram/io_dmi_rd_data[9] ;
input \asic/lsdram/msdram/io_dmi_rd_data[8] ;
input \asic/lsdram/msdram/io_dmi_rd_data[7] ;
input \asic/lsdram/msdram/io_dmi_rd_data[6] ;
input \asic/lsdram/msdram/io_dmi_rd_data[5] ;
input \asic/lsdram/msdram/io_dmi_rd_data[4] ;
input \asic/lsdram/msdram/io_dmi_rd_data[3] ;
input \asic/lsdram/msdram/io_dmi_rd_data[2] ;
input \asic/lsdram/msdram/io_dmi_rd_data[1] ;
input \asic/lsdram/msdram/io_dmi_rd_data[0] ;
input \asic/lsdram/msdram/io_in_rdata_r[255] ;
input \asic/lsdram/msdram/io_in_rdata_r[254] ;
input \asic/lsdram/msdram/io_in_rdata_r[253] ;
input \asic/lsdram/msdram/io_in_rdata_r[252] ;
input \asic/lsdram/msdram/io_in_rdata_r[251] ;
input \asic/lsdram/msdram/io_in_rdata_r[250] ;
input \asic/lsdram/msdram/io_in_rdata_r[249] ;
input \asic/lsdram/msdram/io_in_rdata_r[248] ;
input \asic/lsdram/msdram/io_in_rdata_r[247] ;
input \asic/lsdram/msdram/io_in_rdata_r[246] ;
input \asic/lsdram/msdram/io_in_rdata_r[245] ;
input \asic/lsdram/msdram/io_in_rdata_r[244] ;
input \asic/lsdram/msdram/io_in_rdata_r[243] ;
input \asic/lsdram/msdram/io_in_rdata_r[242] ;
input \asic/lsdram/msdram/io_in_rdata_r[241] ;
input \asic/lsdram/msdram/io_in_rdata_r[240] ;
input \asic/lsdram/msdram/io_in_rdata_r[239] ;
input \asic/lsdram/msdram/io_in_rdata_r[238] ;
input \asic/lsdram/msdram/io_in_rdata_r[237] ;
input \asic/lsdram/msdram/io_in_rdata_r[236] ;
input \asic/lsdram/msdram/io_in_rdata_r[235] ;
input \asic/lsdram/msdram/io_in_rdata_r[234] ;
input \asic/lsdram/msdram/io_in_rdata_r[233] ;
input \asic/lsdram/msdram/io_in_rdata_r[232] ;
input \asic/lsdram/msdram/io_in_rdata_r[231] ;
input \asic/lsdram/msdram/io_in_rdata_r[230] ;
input \asic/lsdram/msdram/io_in_rdata_r[229] ;
input \asic/lsdram/msdram/io_in_rdata_r[228] ;
input \asic/lsdram/msdram/io_in_rdata_r[227] ;
input \asic/lsdram/msdram/io_in_rdata_r[226] ;
input \asic/lsdram/msdram/io_in_rdata_r[225] ;
input \asic/lsdram/msdram/io_in_rdata_r[224] ;
input \asic/lsdram/msdram/io_in_rdata_r[223] ;
input \asic/lsdram/msdram/io_in_rdata_r[222] ;
input \asic/lsdram/msdram/io_in_rdata_r[221] ;
input \asic/lsdram/msdram/io_in_rdata_r[220] ;
input \asic/lsdram/msdram/io_in_rdata_r[219] ;
input \asic/lsdram/msdram/io_in_rdata_r[218] ;
input \asic/lsdram/msdram/io_in_rdata_r[217] ;
input \asic/lsdram/msdram/io_in_rdata_r[216] ;
input \asic/lsdram/msdram/io_in_rdata_r[215] ;
input \asic/lsdram/msdram/io_in_rdata_r[214] ;
input \asic/lsdram/msdram/io_in_rdata_r[213] ;
input \asic/lsdram/msdram/io_in_rdata_r[212] ;
input \asic/lsdram/msdram/io_in_rdata_r[211] ;
input \asic/lsdram/msdram/io_in_rdata_r[210] ;
input \asic/lsdram/msdram/io_in_rdata_r[209] ;
input \asic/lsdram/msdram/io_in_rdata_r[208] ;
input \asic/lsdram/msdram/io_in_rdata_r[207] ;
input \asic/lsdram/msdram/io_in_rdata_r[206] ;
input \asic/lsdram/msdram/io_in_rdata_r[205] ;
input \asic/lsdram/msdram/io_in_rdata_r[204] ;
input \asic/lsdram/msdram/io_in_rdata_r[203] ;
input \asic/lsdram/msdram/io_in_rdata_r[202] ;
input \asic/lsdram/msdram/io_in_rdata_r[201] ;
input \asic/lsdram/msdram/io_in_rdata_r[200] ;
input \asic/lsdram/msdram/io_in_rdata_r[199] ;
input \asic/lsdram/msdram/io_in_rdata_r[198] ;
input \asic/lsdram/msdram/io_in_rdata_r[197] ;
input \asic/lsdram/msdram/io_in_rdata_r[196] ;
input \asic/lsdram/msdram/io_in_rdata_r[195] ;
input \asic/lsdram/msdram/io_in_rdata_r[194] ;
input \asic/lsdram/msdram/io_in_rdata_r[193] ;
input \asic/lsdram/msdram/io_in_rdata_r[192] ;
input \asic/lsdram/msdram/io_in_rdata_r[191] ;
input \asic/lsdram/msdram/io_in_rdata_r[190] ;
input \asic/lsdram/msdram/io_in_rdata_r[189] ;
input \asic/lsdram/msdram/io_in_rdata_r[188] ;
input \asic/lsdram/msdram/io_in_rdata_r[187] ;
input \asic/lsdram/msdram/io_in_rdata_r[186] ;
input \asic/lsdram/msdram/io_in_rdata_r[185] ;
input \asic/lsdram/msdram/io_in_rdata_r[184] ;
input \asic/lsdram/msdram/io_in_rdata_r[183] ;
input \asic/lsdram/msdram/io_in_rdata_r[182] ;
input \asic/lsdram/msdram/io_in_rdata_r[181] ;
input \asic/lsdram/msdram/io_in_rdata_r[180] ;
input \asic/lsdram/msdram/io_in_rdata_r[179] ;
input \asic/lsdram/msdram/io_in_rdata_r[178] ;
input \asic/lsdram/msdram/io_in_rdata_r[177] ;
input \asic/lsdram/msdram/io_in_rdata_r[176] ;
input \asic/lsdram/msdram/io_in_rdata_r[175] ;
input \asic/lsdram/msdram/io_in_rdata_r[174] ;
input \asic/lsdram/msdram/io_in_rdata_r[173] ;
input \asic/lsdram/msdram/io_in_rdata_r[172] ;
input \asic/lsdram/msdram/io_in_rdata_r[171] ;
input \asic/lsdram/msdram/io_in_rdata_r[170] ;
input \asic/lsdram/msdram/io_in_rdata_r[169] ;
input \asic/lsdram/msdram/io_in_rdata_r[168] ;
input \asic/lsdram/msdram/io_in_rdata_r[167] ;
input \asic/lsdram/msdram/io_in_rdata_r[166] ;
input \asic/lsdram/msdram/io_in_rdata_r[165] ;
input \asic/lsdram/msdram/io_in_rdata_r[164] ;
input \asic/lsdram/msdram/io_in_rdata_r[163] ;
input \asic/lsdram/msdram/io_in_rdata_r[162] ;
input \asic/lsdram/msdram/io_in_rdata_r[161] ;
input \asic/lsdram/msdram/io_in_rdata_r[160] ;
input \asic/lsdram/msdram/io_in_rdata_r[159] ;
input \asic/lsdram/msdram/io_in_rdata_r[158] ;
input \asic/lsdram/msdram/io_in_rdata_r[157] ;
input \asic/lsdram/msdram/io_in_rdata_r[156] ;
input \asic/lsdram/msdram/io_in_rdata_r[155] ;
input \asic/lsdram/msdram/io_in_rdata_r[154] ;
input \asic/lsdram/msdram/io_in_rdata_r[153] ;
input \asic/lsdram/msdram/io_in_rdata_r[152] ;
input \asic/lsdram/msdram/io_in_rdata_r[151] ;
input \asic/lsdram/msdram/io_in_rdata_r[150] ;
input \asic/lsdram/msdram/io_in_rdata_r[149] ;
input \asic/lsdram/msdram/io_in_rdata_r[148] ;
input \asic/lsdram/msdram/io_in_rdata_r[147] ;
input \asic/lsdram/msdram/io_in_rdata_r[146] ;
input \asic/lsdram/msdram/io_in_rdata_r[145] ;
input \asic/lsdram/msdram/io_in_rdata_r[144] ;
input \asic/lsdram/msdram/io_in_rdata_r[143] ;
input \asic/lsdram/msdram/io_in_rdata_r[142] ;
input \asic/lsdram/msdram/io_in_rdata_r[141] ;
input \asic/lsdram/msdram/io_in_rdata_r[140] ;
input \asic/lsdram/msdram/io_in_rdata_r[139] ;
input \asic/lsdram/msdram/io_in_rdata_r[138] ;
input \asic/lsdram/msdram/io_in_rdata_r[137] ;
input \asic/lsdram/msdram/io_in_rdata_r[136] ;
input \asic/lsdram/msdram/io_in_rdata_r[135] ;
input \asic/lsdram/msdram/io_in_rdata_r[134] ;
input \asic/lsdram/msdram/io_in_rdata_r[133] ;
input \asic/lsdram/msdram/io_in_rdata_r[132] ;
input \asic/lsdram/msdram/io_in_rdata_r[131] ;
input \asic/lsdram/msdram/io_in_rdata_r[130] ;
input \asic/lsdram/msdram/io_in_rdata_r[129] ;
input \asic/lsdram/msdram/io_in_rdata_r[128] ;
input \asic/lsdram/msdram/io_in_rdata_r[127] ;
input \asic/lsdram/msdram/io_in_rdata_r[126] ;
input \asic/lsdram/msdram/io_in_rdata_r[125] ;
input \asic/lsdram/msdram/io_in_rdata_r[124] ;
input \asic/lsdram/msdram/io_in_rdata_r[123] ;
input \asic/lsdram/msdram/io_in_rdata_r[122] ;
input \asic/lsdram/msdram/io_in_rdata_r[121] ;
input \asic/lsdram/msdram/io_in_rdata_r[120] ;
input \asic/lsdram/msdram/io_in_rdata_r[119] ;
input \asic/lsdram/msdram/io_in_rdata_r[118] ;
input \asic/lsdram/msdram/io_in_rdata_r[117] ;
input \asic/lsdram/msdram/io_in_rdata_r[116] ;
input \asic/lsdram/msdram/io_in_rdata_r[115] ;
input \asic/lsdram/msdram/io_in_rdata_r[114] ;
input \asic/lsdram/msdram/io_in_rdata_r[113] ;
input \asic/lsdram/msdram/io_in_rdata_r[112] ;
input \asic/lsdram/msdram/io_in_rdata_r[111] ;
input \asic/lsdram/msdram/io_in_rdata_r[110] ;
input \asic/lsdram/msdram/io_in_rdata_r[109] ;
input \asic/lsdram/msdram/io_in_rdata_r[108] ;
input \asic/lsdram/msdram/io_in_rdata_r[107] ;
input \asic/lsdram/msdram/io_in_rdata_r[106] ;
input \asic/lsdram/msdram/io_in_rdata_r[105] ;
input \asic/lsdram/msdram/io_in_rdata_r[104] ;
input \asic/lsdram/msdram/io_in_rdata_r[103] ;
input \asic/lsdram/msdram/io_in_rdata_r[102] ;
input \asic/lsdram/msdram/io_in_rdata_r[101] ;
input \asic/lsdram/msdram/io_in_rdata_r[100] ;
input \asic/lsdram/msdram/io_in_rdata_r[99] ;
input \asic/lsdram/msdram/io_in_rdata_r[98] ;
input \asic/lsdram/msdram/io_in_rdata_r[97] ;
input \asic/lsdram/msdram/io_in_rdata_r[96] ;
input \asic/lsdram/msdram/io_in_rdata_r[95] ;
input \asic/lsdram/msdram/io_in_rdata_r[94] ;
input \asic/lsdram/msdram/io_in_rdata_r[93] ;
input \asic/lsdram/msdram/io_in_rdata_r[92] ;
input \asic/lsdram/msdram/io_in_rdata_r[91] ;
input \asic/lsdram/msdram/io_in_rdata_r[90] ;
input \asic/lsdram/msdram/io_in_rdata_r[89] ;
input \asic/lsdram/msdram/io_in_rdata_r[88] ;
input \asic/lsdram/msdram/io_in_rdata_r[87] ;
input \asic/lsdram/msdram/io_in_rdata_r[86] ;
input \asic/lsdram/msdram/io_in_rdata_r[85] ;
input \asic/lsdram/msdram/io_in_rdata_r[84] ;
input \asic/lsdram/msdram/io_in_rdata_r[83] ;
input \asic/lsdram/msdram/io_in_rdata_r[82] ;
input \asic/lsdram/msdram/io_in_rdata_r[81] ;
input \asic/lsdram/msdram/io_in_rdata_r[80] ;
input \asic/lsdram/msdram/io_in_rdata_r[79] ;
input \asic/lsdram/msdram/io_in_rdata_r[78] ;
input \asic/lsdram/msdram/io_in_rdata_r[77] ;
input \asic/lsdram/msdram/io_in_rdata_r[76] ;
input \asic/lsdram/msdram/io_in_rdata_r[75] ;
input \asic/lsdram/msdram/io_in_rdata_r[74] ;
input \asic/lsdram/msdram/io_in_rdata_r[73] ;
input \asic/lsdram/msdram/io_in_rdata_r[72] ;
input \asic/lsdram/msdram/io_in_rdata_r[71] ;
input \asic/lsdram/msdram/io_in_rdata_r[70] ;
input \asic/lsdram/msdram/io_in_rdata_r[69] ;
input \asic/lsdram/msdram/io_in_rdata_r[68] ;
input \asic/lsdram/msdram/io_in_rdata_r[67] ;
input \asic/lsdram/msdram/io_in_rdata_r[66] ;
input \asic/lsdram/msdram/io_in_rdata_r[65] ;
input \asic/lsdram/msdram/io_in_rdata_r[64] ;
input \asic/lsdram/msdram/io_in_rdata_r[63] ;
input \asic/lsdram/msdram/io_in_rdata_r[62] ;
input \asic/lsdram/msdram/io_in_rdata_r[61] ;
input \asic/lsdram/msdram/io_in_rdata_r[60] ;
input \asic/lsdram/msdram/io_in_rdata_r[59] ;
input \asic/lsdram/msdram/io_in_rdata_r[58] ;
input \asic/lsdram/msdram/io_in_rdata_r[57] ;
input \asic/lsdram/msdram/io_in_rdata_r[56] ;
input \asic/lsdram/msdram/io_in_rdata_r[55] ;
input \asic/lsdram/msdram/io_in_rdata_r[54] ;
input \asic/lsdram/msdram/io_in_rdata_r[53] ;
input \asic/lsdram/msdram/io_in_rdata_r[52] ;
input \asic/lsdram/msdram/io_in_rdata_r[51] ;
input \asic/lsdram/msdram/io_in_rdata_r[50] ;
input \asic/lsdram/msdram/io_in_rdata_r[49] ;
input \asic/lsdram/msdram/io_in_rdata_r[48] ;
input \asic/lsdram/msdram/io_in_rdata_r[47] ;
input \asic/lsdram/msdram/io_in_rdata_r[46] ;
input \asic/lsdram/msdram/io_in_rdata_r[45] ;
input \asic/lsdram/msdram/io_in_rdata_r[44] ;
input \asic/lsdram/msdram/io_in_rdata_r[43] ;
input \asic/lsdram/msdram/io_in_rdata_r[42] ;
input \asic/lsdram/msdram/io_in_rdata_r[41] ;
input \asic/lsdram/msdram/io_in_rdata_r[40] ;
input \asic/lsdram/msdram/io_in_rdata_r[39] ;
input \asic/lsdram/msdram/io_in_rdata_r[38] ;
input \asic/lsdram/msdram/io_in_rdata_r[37] ;
input \asic/lsdram/msdram/io_in_rdata_r[36] ;
input \asic/lsdram/msdram/io_in_rdata_r[35] ;
input \asic/lsdram/msdram/io_in_rdata_r[34] ;
input \asic/lsdram/msdram/io_in_rdata_r[33] ;
input \asic/lsdram/msdram/io_in_rdata_r[32] ;
input \asic/lsdram/msdram/io_in_rdata_r[31] ;
input \asic/lsdram/msdram/io_in_rdata_r[30] ;
input \asic/lsdram/msdram/io_in_rdata_r[29] ;
input \asic/lsdram/msdram/io_in_rdata_r[28] ;
input \asic/lsdram/msdram/io_in_rdata_r[27] ;
input \asic/lsdram/msdram/io_in_rdata_r[26] ;
input \asic/lsdram/msdram/io_in_rdata_r[25] ;
input \asic/lsdram/msdram/io_in_rdata_r[24] ;
input \asic/lsdram/msdram/io_in_rdata_r[23] ;
input \asic/lsdram/msdram/io_in_rdata_r[22] ;
input \asic/lsdram/msdram/io_in_rdata_r[21] ;
input \asic/lsdram/msdram/io_in_rdata_r[20] ;
input \asic/lsdram/msdram/io_in_rdata_r[19] ;
input \asic/lsdram/msdram/io_in_rdata_r[18] ;
input \asic/lsdram/msdram/io_in_rdata_r[17] ;
input \asic/lsdram/msdram/io_in_rdata_r[16] ;
input \asic/lsdram/msdram/io_in_rdata_r[15] ;
input \asic/lsdram/msdram/io_in_rdata_r[14] ;
input \asic/lsdram/msdram/io_in_rdata_r[13] ;
input \asic/lsdram/msdram/io_in_rdata_r[12] ;
input \asic/lsdram/msdram/io_in_rdata_r[11] ;
input \asic/lsdram/msdram/io_in_rdata_r[10] ;
input \asic/lsdram/msdram/io_in_rdata_r[9] ;
input \asic/lsdram/msdram/io_in_rdata_r[8] ;
input \asic/lsdram/msdram/io_in_rdata_r[7] ;
input \asic/lsdram/msdram/io_in_rdata_r[6] ;
input \asic/lsdram/msdram/io_in_rdata_r[5] ;
input \asic/lsdram/msdram/io_in_rdata_r[4] ;
input \asic/lsdram/msdram/io_in_rdata_r[3] ;
input \asic/lsdram/msdram/io_in_rdata_r[2] ;
input \asic/lsdram/msdram/io_in_rdata_r[1] ;
input \asic/lsdram/msdram/io_in_rdata_r[0] ;
input \asic/lsdram/msdram/io_clk_out ;
input \asic/lsdram/msdram/io_in_awready ;
input \asic/lsdram/msdram/io_in_awvalid ;
input \asic/lsdram/msdram/io_in_wready ;
input \asic/lsdram/msdram/io_in_wvalid ;
input \asic/lsdram/msdram/io_in_bready ;
input \asic/lsdram/msdram/io_in_bvalid ;
input \asic/lsdram/msdram/io_in_arready ;
input \asic/lsdram/msdram/io_in_arvalid ;
input \asic/lsdram/msdram/io_in_rready ;
input \asic/lsdram/msdram/io_in_rvalid ;
input \asic/lsdram/msdram/io_dmi_cmd_en ;
input \asic/lsdram/msdram/io_dmi_wr_data_en ;
input \asic/lsdram/msdram/io_dmi_wr_data_end ;
input \asic/lsdram/msdram/io_dmi_clk_out ;
input \asic/lsdram/msdram/io_dmi_init_calib_complete ;
input \asic/lsdram/msdram/io_dmi_cmd_ready ;
input \asic/lsdram/msdram/io_dmi_wr_data_rdy ;
input \asic/lsdram/msdram/io_dmi_rd_data_valid ;
input clock;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \asic/cpu/cpu/if_stage/fs_pc[31] ;
wire \asic/cpu/cpu/if_stage/fs_pc[30] ;
wire \asic/cpu/cpu/if_stage/fs_pc[29] ;
wire \asic/cpu/cpu/if_stage/fs_pc[28] ;
wire \asic/cpu/cpu/if_stage/fs_pc[27] ;
wire \asic/cpu/cpu/if_stage/fs_pc[26] ;
wire \asic/cpu/cpu/if_stage/fs_pc[25] ;
wire \asic/cpu/cpu/if_stage/fs_pc[24] ;
wire \asic/cpu/cpu/if_stage/fs_pc[23] ;
wire \asic/cpu/cpu/if_stage/fs_pc[22] ;
wire \asic/cpu/cpu/if_stage/fs_pc[21] ;
wire \asic/cpu/cpu/if_stage/fs_pc[20] ;
wire \asic/cpu/cpu/if_stage/fs_pc[19] ;
wire \asic/cpu/cpu/if_stage/fs_pc[18] ;
wire \asic/cpu/cpu/if_stage/fs_pc[17] ;
wire \asic/cpu/cpu/if_stage/fs_pc[16] ;
wire \asic/cpu/cpu/if_stage/fs_pc[15] ;
wire \asic/cpu/cpu/if_stage/fs_pc[14] ;
wire \asic/cpu/cpu/if_stage/fs_pc[13] ;
wire \asic/cpu/cpu/if_stage/fs_pc[12] ;
wire \asic/cpu/cpu/if_stage/fs_pc[11] ;
wire \asic/cpu/cpu/if_stage/fs_pc[10] ;
wire \asic/cpu/cpu/if_stage/fs_pc[9] ;
wire \asic/cpu/cpu/if_stage/fs_pc[8] ;
wire \asic/cpu/cpu/if_stage/fs_pc[7] ;
wire \asic/cpu/cpu/if_stage/fs_pc[6] ;
wire \asic/cpu/cpu/if_stage/fs_pc[5] ;
wire \asic/cpu/cpu/if_stage/fs_pc[4] ;
wire \asic/cpu/cpu/if_stage/fs_pc[3] ;
wire \asic/cpu/cpu/if_stage/fs_pc[2] ;
wire \asic/cpu/cpu/if_stage/fs_pc[1] ;
wire \asic/cpu/cpu/if_stage/fs_pc[0] ;
wire \asic/cpu/cpu/if_stage/fs_inst[31] ;
wire \asic/cpu/cpu/if_stage/fs_inst[30] ;
wire \asic/cpu/cpu/if_stage/fs_inst[29] ;
wire \asic/cpu/cpu/if_stage/fs_inst[28] ;
wire \asic/cpu/cpu/if_stage/fs_inst[27] ;
wire \asic/cpu/cpu/if_stage/fs_inst[26] ;
wire \asic/cpu/cpu/if_stage/fs_inst[25] ;
wire \asic/cpu/cpu/if_stage/fs_inst[24] ;
wire \asic/cpu/cpu/if_stage/fs_inst[23] ;
wire \asic/cpu/cpu/if_stage/fs_inst[22] ;
wire \asic/cpu/cpu/if_stage/fs_inst[21] ;
wire \asic/cpu/cpu/if_stage/fs_inst[20] ;
wire \asic/cpu/cpu/if_stage/fs_inst[19] ;
wire \asic/cpu/cpu/if_stage/fs_inst[18] ;
wire \asic/cpu/cpu/if_stage/fs_inst[17] ;
wire \asic/cpu/cpu/if_stage/fs_inst[16] ;
wire \asic/cpu/cpu/if_stage/fs_inst[15] ;
wire \asic/cpu/cpu/if_stage/fs_inst[14] ;
wire \asic/cpu/cpu/if_stage/fs_inst[13] ;
wire \asic/cpu/cpu/if_stage/fs_inst[12] ;
wire \asic/cpu/cpu/if_stage/fs_inst[11] ;
wire \asic/cpu/cpu/if_stage/fs_inst[10] ;
wire \asic/cpu/cpu/if_stage/fs_inst[9] ;
wire \asic/cpu/cpu/if_stage/fs_inst[8] ;
wire \asic/cpu/cpu/if_stage/fs_inst[7] ;
wire \asic/cpu/cpu/if_stage/fs_inst[6] ;
wire \asic/cpu/cpu/if_stage/fs_inst[5] ;
wire \asic/cpu/cpu/if_stage/fs_inst[4] ;
wire \asic/cpu/cpu/if_stage/fs_inst[3] ;
wire \asic/cpu/cpu/if_stage/fs_inst[2] ;
wire \asic/cpu/cpu/if_stage/fs_inst[1] ;
wire \asic/cpu/cpu/if_stage/fs_inst[0] ;
wire \asic/lsdram/msdram/io_in_awid[3] ;
wire \asic/lsdram/msdram/io_in_awid[2] ;
wire \asic/lsdram/msdram/io_in_awid[1] ;
wire \asic/lsdram/msdram/io_in_awid[0] ;
wire \asic/lsdram/msdram/io_in_awaddr[31] ;
wire \asic/lsdram/msdram/io_in_awaddr[30] ;
wire \asic/lsdram/msdram/io_in_awaddr[29] ;
wire \asic/lsdram/msdram/io_in_awaddr[28] ;
wire \asic/lsdram/msdram/io_in_awaddr[27] ;
wire \asic/lsdram/msdram/io_in_awaddr[26] ;
wire \asic/lsdram/msdram/io_in_awaddr[25] ;
wire \asic/lsdram/msdram/io_in_awaddr[24] ;
wire \asic/lsdram/msdram/io_in_awaddr[23] ;
wire \asic/lsdram/msdram/io_in_awaddr[22] ;
wire \asic/lsdram/msdram/io_in_awaddr[21] ;
wire \asic/lsdram/msdram/io_in_awaddr[20] ;
wire \asic/lsdram/msdram/io_in_awaddr[19] ;
wire \asic/lsdram/msdram/io_in_awaddr[18] ;
wire \asic/lsdram/msdram/io_in_awaddr[17] ;
wire \asic/lsdram/msdram/io_in_awaddr[16] ;
wire \asic/lsdram/msdram/io_in_awaddr[15] ;
wire \asic/lsdram/msdram/io_in_awaddr[14] ;
wire \asic/lsdram/msdram/io_in_awaddr[13] ;
wire \asic/lsdram/msdram/io_in_awaddr[12] ;
wire \asic/lsdram/msdram/io_in_awaddr[11] ;
wire \asic/lsdram/msdram/io_in_awaddr[10] ;
wire \asic/lsdram/msdram/io_in_awaddr[9] ;
wire \asic/lsdram/msdram/io_in_awaddr[8] ;
wire \asic/lsdram/msdram/io_in_awaddr[7] ;
wire \asic/lsdram/msdram/io_in_awaddr[6] ;
wire \asic/lsdram/msdram/io_in_awaddr[5] ;
wire \asic/lsdram/msdram/io_in_awaddr[4] ;
wire \asic/lsdram/msdram/io_in_awaddr[3] ;
wire \asic/lsdram/msdram/io_in_awaddr[2] ;
wire \asic/lsdram/msdram/io_in_awaddr[1] ;
wire \asic/lsdram/msdram/io_in_awaddr[0] ;
wire \asic/lsdram/msdram/io_in_awlen[7] ;
wire \asic/lsdram/msdram/io_in_awlen[6] ;
wire \asic/lsdram/msdram/io_in_awlen[5] ;
wire \asic/lsdram/msdram/io_in_awlen[4] ;
wire \asic/lsdram/msdram/io_in_awlen[3] ;
wire \asic/lsdram/msdram/io_in_awlen[2] ;
wire \asic/lsdram/msdram/io_in_awlen[1] ;
wire \asic/lsdram/msdram/io_in_awlen[0] ;
wire \asic/lsdram/msdram/io_in_awsize[2] ;
wire \asic/lsdram/msdram/io_in_awsize[1] ;
wire \asic/lsdram/msdram/io_in_awsize[0] ;
wire \asic/lsdram/msdram/io_in_wdata[31] ;
wire \asic/lsdram/msdram/io_in_wdata[30] ;
wire \asic/lsdram/msdram/io_in_wdata[29] ;
wire \asic/lsdram/msdram/io_in_wdata[28] ;
wire \asic/lsdram/msdram/io_in_wdata[27] ;
wire \asic/lsdram/msdram/io_in_wdata[26] ;
wire \asic/lsdram/msdram/io_in_wdata[25] ;
wire \asic/lsdram/msdram/io_in_wdata[24] ;
wire \asic/lsdram/msdram/io_in_wdata[23] ;
wire \asic/lsdram/msdram/io_in_wdata[22] ;
wire \asic/lsdram/msdram/io_in_wdata[21] ;
wire \asic/lsdram/msdram/io_in_wdata[20] ;
wire \asic/lsdram/msdram/io_in_wdata[19] ;
wire \asic/lsdram/msdram/io_in_wdata[18] ;
wire \asic/lsdram/msdram/io_in_wdata[17] ;
wire \asic/lsdram/msdram/io_in_wdata[16] ;
wire \asic/lsdram/msdram/io_in_wdata[15] ;
wire \asic/lsdram/msdram/io_in_wdata[14] ;
wire \asic/lsdram/msdram/io_in_wdata[13] ;
wire \asic/lsdram/msdram/io_in_wdata[12] ;
wire \asic/lsdram/msdram/io_in_wdata[11] ;
wire \asic/lsdram/msdram/io_in_wdata[10] ;
wire \asic/lsdram/msdram/io_in_wdata[9] ;
wire \asic/lsdram/msdram/io_in_wdata[8] ;
wire \asic/lsdram/msdram/io_in_wdata[7] ;
wire \asic/lsdram/msdram/io_in_wdata[6] ;
wire \asic/lsdram/msdram/io_in_wdata[5] ;
wire \asic/lsdram/msdram/io_in_wdata[4] ;
wire \asic/lsdram/msdram/io_in_wdata[3] ;
wire \asic/lsdram/msdram/io_in_wdata[2] ;
wire \asic/lsdram/msdram/io_in_wdata[1] ;
wire \asic/lsdram/msdram/io_in_wdata[0] ;
wire \asic/lsdram/msdram/io_in_wstrb[3] ;
wire \asic/lsdram/msdram/io_in_wstrb[2] ;
wire \asic/lsdram/msdram/io_in_wstrb[1] ;
wire \asic/lsdram/msdram/io_in_wstrb[0] ;
wire \asic/lsdram/msdram/io_in_bid[3] ;
wire \asic/lsdram/msdram/io_in_bid[2] ;
wire \asic/lsdram/msdram/io_in_bid[1] ;
wire \asic/lsdram/msdram/io_in_bid[0] ;
wire \asic/lsdram/msdram/io_in_arid[3] ;
wire \asic/lsdram/msdram/io_in_arid[2] ;
wire \asic/lsdram/msdram/io_in_arid[1] ;
wire \asic/lsdram/msdram/io_in_arid[0] ;
wire \asic/lsdram/msdram/io_in_araddr[31] ;
wire \asic/lsdram/msdram/io_in_araddr[30] ;
wire \asic/lsdram/msdram/io_in_araddr[29] ;
wire \asic/lsdram/msdram/io_in_araddr[28] ;
wire \asic/lsdram/msdram/io_in_araddr[27] ;
wire \asic/lsdram/msdram/io_in_araddr[26] ;
wire \asic/lsdram/msdram/io_in_araddr[25] ;
wire \asic/lsdram/msdram/io_in_araddr[24] ;
wire \asic/lsdram/msdram/io_in_araddr[23] ;
wire \asic/lsdram/msdram/io_in_araddr[22] ;
wire \asic/lsdram/msdram/io_in_araddr[21] ;
wire \asic/lsdram/msdram/io_in_araddr[20] ;
wire \asic/lsdram/msdram/io_in_araddr[19] ;
wire \asic/lsdram/msdram/io_in_araddr[18] ;
wire \asic/lsdram/msdram/io_in_araddr[17] ;
wire \asic/lsdram/msdram/io_in_araddr[16] ;
wire \asic/lsdram/msdram/io_in_araddr[15] ;
wire \asic/lsdram/msdram/io_in_araddr[14] ;
wire \asic/lsdram/msdram/io_in_araddr[13] ;
wire \asic/lsdram/msdram/io_in_araddr[12] ;
wire \asic/lsdram/msdram/io_in_araddr[11] ;
wire \asic/lsdram/msdram/io_in_araddr[10] ;
wire \asic/lsdram/msdram/io_in_araddr[9] ;
wire \asic/lsdram/msdram/io_in_araddr[8] ;
wire \asic/lsdram/msdram/io_in_araddr[7] ;
wire \asic/lsdram/msdram/io_in_araddr[6] ;
wire \asic/lsdram/msdram/io_in_araddr[5] ;
wire \asic/lsdram/msdram/io_in_araddr[4] ;
wire \asic/lsdram/msdram/io_in_araddr[3] ;
wire \asic/lsdram/msdram/io_in_araddr[2] ;
wire \asic/lsdram/msdram/io_in_araddr[1] ;
wire \asic/lsdram/msdram/io_in_araddr[0] ;
wire \asic/lsdram/msdram/io_in_arlen[7] ;
wire \asic/lsdram/msdram/io_in_arlen[6] ;
wire \asic/lsdram/msdram/io_in_arlen[5] ;
wire \asic/lsdram/msdram/io_in_arlen[4] ;
wire \asic/lsdram/msdram/io_in_arlen[3] ;
wire \asic/lsdram/msdram/io_in_arlen[2] ;
wire \asic/lsdram/msdram/io_in_arlen[1] ;
wire \asic/lsdram/msdram/io_in_arlen[0] ;
wire \asic/lsdram/msdram/io_in_arsize[2] ;
wire \asic/lsdram/msdram/io_in_arsize[1] ;
wire \asic/lsdram/msdram/io_in_arsize[0] ;
wire \asic/lsdram/msdram/io_in_rid[3] ;
wire \asic/lsdram/msdram/io_in_rid[2] ;
wire \asic/lsdram/msdram/io_in_rid[1] ;
wire \asic/lsdram/msdram/io_in_rid[0] ;
wire \asic/lsdram/msdram/io_in_rdata[31] ;
wire \asic/lsdram/msdram/io_in_rdata[30] ;
wire \asic/lsdram/msdram/io_in_rdata[29] ;
wire \asic/lsdram/msdram/io_in_rdata[28] ;
wire \asic/lsdram/msdram/io_in_rdata[27] ;
wire \asic/lsdram/msdram/io_in_rdata[26] ;
wire \asic/lsdram/msdram/io_in_rdata[25] ;
wire \asic/lsdram/msdram/io_in_rdata[24] ;
wire \asic/lsdram/msdram/io_in_rdata[23] ;
wire \asic/lsdram/msdram/io_in_rdata[22] ;
wire \asic/lsdram/msdram/io_in_rdata[21] ;
wire \asic/lsdram/msdram/io_in_rdata[20] ;
wire \asic/lsdram/msdram/io_in_rdata[19] ;
wire \asic/lsdram/msdram/io_in_rdata[18] ;
wire \asic/lsdram/msdram/io_in_rdata[17] ;
wire \asic/lsdram/msdram/io_in_rdata[16] ;
wire \asic/lsdram/msdram/io_in_rdata[15] ;
wire \asic/lsdram/msdram/io_in_rdata[14] ;
wire \asic/lsdram/msdram/io_in_rdata[13] ;
wire \asic/lsdram/msdram/io_in_rdata[12] ;
wire \asic/lsdram/msdram/io_in_rdata[11] ;
wire \asic/lsdram/msdram/io_in_rdata[10] ;
wire \asic/lsdram/msdram/io_in_rdata[9] ;
wire \asic/lsdram/msdram/io_in_rdata[8] ;
wire \asic/lsdram/msdram/io_in_rdata[7] ;
wire \asic/lsdram/msdram/io_in_rdata[6] ;
wire \asic/lsdram/msdram/io_in_rdata[5] ;
wire \asic/lsdram/msdram/io_in_rdata[4] ;
wire \asic/lsdram/msdram/io_in_rdata[3] ;
wire \asic/lsdram/msdram/io_in_rdata[2] ;
wire \asic/lsdram/msdram/io_in_rdata[1] ;
wire \asic/lsdram/msdram/io_in_rdata[0] ;
wire \asic/lsdram/msdram/io_dmi_cmd[2] ;
wire \asic/lsdram/msdram/io_dmi_cmd[1] ;
wire \asic/lsdram/msdram/io_dmi_cmd[0] ;
wire \asic/lsdram/msdram/io_dmi_addr[28] ;
wire \asic/lsdram/msdram/io_dmi_addr[27] ;
wire \asic/lsdram/msdram/io_dmi_addr[26] ;
wire \asic/lsdram/msdram/io_dmi_addr[25] ;
wire \asic/lsdram/msdram/io_dmi_addr[24] ;
wire \asic/lsdram/msdram/io_dmi_addr[23] ;
wire \asic/lsdram/msdram/io_dmi_addr[22] ;
wire \asic/lsdram/msdram/io_dmi_addr[21] ;
wire \asic/lsdram/msdram/io_dmi_addr[20] ;
wire \asic/lsdram/msdram/io_dmi_addr[19] ;
wire \asic/lsdram/msdram/io_dmi_addr[18] ;
wire \asic/lsdram/msdram/io_dmi_addr[17] ;
wire \asic/lsdram/msdram/io_dmi_addr[16] ;
wire \asic/lsdram/msdram/io_dmi_addr[15] ;
wire \asic/lsdram/msdram/io_dmi_addr[14] ;
wire \asic/lsdram/msdram/io_dmi_addr[13] ;
wire \asic/lsdram/msdram/io_dmi_addr[12] ;
wire \asic/lsdram/msdram/io_dmi_addr[11] ;
wire \asic/lsdram/msdram/io_dmi_addr[10] ;
wire \asic/lsdram/msdram/io_dmi_addr[9] ;
wire \asic/lsdram/msdram/io_dmi_addr[8] ;
wire \asic/lsdram/msdram/io_dmi_addr[7] ;
wire \asic/lsdram/msdram/io_dmi_addr[6] ;
wire \asic/lsdram/msdram/io_dmi_addr[5] ;
wire \asic/lsdram/msdram/io_dmi_addr[4] ;
wire \asic/lsdram/msdram/io_dmi_addr[3] ;
wire \asic/lsdram/msdram/io_dmi_addr[2] ;
wire \asic/lsdram/msdram/io_dmi_addr[1] ;
wire \asic/lsdram/msdram/io_dmi_addr[0] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[255] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[254] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[253] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[252] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[251] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[250] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[249] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[248] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[247] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[246] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[245] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[244] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[243] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[242] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[241] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[240] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[239] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[238] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[237] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[236] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[235] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[234] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[233] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[232] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[231] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[230] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[229] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[228] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[227] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[226] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[225] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[224] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[223] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[222] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[221] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[220] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[219] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[218] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[217] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[216] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[215] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[214] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[213] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[212] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[211] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[210] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[209] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[208] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[207] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[206] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[205] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[204] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[203] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[202] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[201] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[200] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[199] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[198] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[197] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[196] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[195] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[194] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[193] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[192] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[191] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[190] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[189] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[188] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[187] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[186] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[185] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[184] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[183] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[182] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[181] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[180] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[179] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[178] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[177] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[176] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[175] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[174] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[173] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[172] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[171] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[170] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[169] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[168] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[167] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[166] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[165] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[164] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[163] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[162] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[161] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[160] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[159] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[158] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[157] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[156] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[155] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[154] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[153] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[152] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[151] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[150] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[149] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[148] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[147] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[146] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[145] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[144] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[143] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[142] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[141] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[140] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[139] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[138] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[137] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[136] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[135] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[134] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[133] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[132] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[131] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[130] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[129] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[128] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[127] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[126] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[125] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[124] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[123] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[122] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[121] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[120] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[119] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[118] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[117] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[116] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[115] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[114] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[113] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[112] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[111] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[110] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[109] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[108] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[107] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[106] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[105] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[104] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[103] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[102] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[101] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[100] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[99] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[98] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[97] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[96] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[95] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[94] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[93] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[92] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[91] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[90] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[89] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[88] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[87] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[86] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[85] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[84] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[83] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[82] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[81] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[80] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[79] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[78] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[77] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[76] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[75] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[74] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[73] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[72] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[71] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[70] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[69] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[68] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[67] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[66] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[65] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[64] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[63] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[62] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[61] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[60] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[59] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[58] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[57] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[56] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[55] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[54] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[53] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[52] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[51] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[50] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[49] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[48] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[47] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[46] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[45] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[44] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[43] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[42] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[41] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[40] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[39] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[38] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[37] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[36] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[35] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[34] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[33] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[32] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[31] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[30] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[29] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[28] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[27] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[26] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[25] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[24] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[23] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[22] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[21] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[20] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[19] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[18] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[17] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[16] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[15] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[14] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[13] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[12] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[11] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[10] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[9] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[8] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[7] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[6] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[5] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[4] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[3] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[2] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[1] ;
wire \asic/lsdram/msdram/io_dmi_wr_data[0] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[31] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[30] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[29] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[28] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[27] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[26] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[25] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[24] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[23] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[22] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[21] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[20] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[19] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[18] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[17] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[16] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[15] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[14] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[13] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[12] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[11] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[10] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[9] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[8] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[7] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[6] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[5] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[4] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[3] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[2] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[1] ;
wire \asic/lsdram/msdram/io_dmi_wr_data_mask[0] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[255] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[254] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[253] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[252] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[251] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[250] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[249] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[248] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[247] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[246] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[245] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[244] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[243] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[242] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[241] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[240] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[239] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[238] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[237] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[236] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[235] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[234] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[233] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[232] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[231] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[230] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[229] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[228] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[227] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[226] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[225] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[224] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[223] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[222] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[221] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[220] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[219] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[218] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[217] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[216] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[215] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[214] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[213] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[212] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[211] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[210] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[209] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[208] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[207] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[206] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[205] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[204] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[203] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[202] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[201] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[200] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[199] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[198] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[197] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[196] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[195] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[194] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[193] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[192] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[191] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[190] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[189] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[188] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[187] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[186] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[185] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[184] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[183] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[182] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[181] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[180] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[179] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[178] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[177] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[176] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[175] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[174] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[173] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[172] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[171] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[170] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[169] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[168] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[167] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[166] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[165] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[164] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[163] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[162] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[161] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[160] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[159] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[158] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[157] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[156] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[155] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[154] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[153] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[152] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[151] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[150] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[149] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[148] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[147] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[146] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[145] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[144] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[143] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[142] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[141] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[140] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[139] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[138] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[137] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[136] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[135] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[134] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[133] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[132] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[131] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[130] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[129] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[128] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[127] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[126] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[125] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[124] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[123] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[122] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[121] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[120] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[119] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[118] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[117] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[116] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[115] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[114] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[113] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[112] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[111] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[110] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[109] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[108] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[107] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[106] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[105] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[104] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[103] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[102] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[101] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[100] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[99] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[98] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[97] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[96] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[95] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[94] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[93] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[92] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[91] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[90] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[89] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[88] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[87] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[86] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[85] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[84] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[83] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[82] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[81] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[80] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[79] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[78] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[77] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[76] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[75] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[74] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[73] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[72] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[71] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[70] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[69] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[68] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[67] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[66] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[65] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[64] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[63] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[62] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[61] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[60] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[59] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[58] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[57] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[56] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[55] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[54] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[53] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[52] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[51] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[50] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[49] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[48] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[47] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[46] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[45] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[44] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[43] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[42] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[41] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[40] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[39] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[38] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[37] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[36] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[35] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[34] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[33] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[32] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[31] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[30] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[29] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[28] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[27] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[26] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[25] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[24] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[23] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[22] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[21] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[20] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[19] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[18] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[17] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[16] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[15] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[14] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[13] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[12] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[11] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[10] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[9] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[8] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[7] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[6] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[5] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[4] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[3] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[2] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[1] ;
wire \asic/lsdram/msdram/io_dmi_rd_data[0] ;
wire \asic/lsdram/msdram/io_in_rdata_r[255] ;
wire \asic/lsdram/msdram/io_in_rdata_r[254] ;
wire \asic/lsdram/msdram/io_in_rdata_r[253] ;
wire \asic/lsdram/msdram/io_in_rdata_r[252] ;
wire \asic/lsdram/msdram/io_in_rdata_r[251] ;
wire \asic/lsdram/msdram/io_in_rdata_r[250] ;
wire \asic/lsdram/msdram/io_in_rdata_r[249] ;
wire \asic/lsdram/msdram/io_in_rdata_r[248] ;
wire \asic/lsdram/msdram/io_in_rdata_r[247] ;
wire \asic/lsdram/msdram/io_in_rdata_r[246] ;
wire \asic/lsdram/msdram/io_in_rdata_r[245] ;
wire \asic/lsdram/msdram/io_in_rdata_r[244] ;
wire \asic/lsdram/msdram/io_in_rdata_r[243] ;
wire \asic/lsdram/msdram/io_in_rdata_r[242] ;
wire \asic/lsdram/msdram/io_in_rdata_r[241] ;
wire \asic/lsdram/msdram/io_in_rdata_r[240] ;
wire \asic/lsdram/msdram/io_in_rdata_r[239] ;
wire \asic/lsdram/msdram/io_in_rdata_r[238] ;
wire \asic/lsdram/msdram/io_in_rdata_r[237] ;
wire \asic/lsdram/msdram/io_in_rdata_r[236] ;
wire \asic/lsdram/msdram/io_in_rdata_r[235] ;
wire \asic/lsdram/msdram/io_in_rdata_r[234] ;
wire \asic/lsdram/msdram/io_in_rdata_r[233] ;
wire \asic/lsdram/msdram/io_in_rdata_r[232] ;
wire \asic/lsdram/msdram/io_in_rdata_r[231] ;
wire \asic/lsdram/msdram/io_in_rdata_r[230] ;
wire \asic/lsdram/msdram/io_in_rdata_r[229] ;
wire \asic/lsdram/msdram/io_in_rdata_r[228] ;
wire \asic/lsdram/msdram/io_in_rdata_r[227] ;
wire \asic/lsdram/msdram/io_in_rdata_r[226] ;
wire \asic/lsdram/msdram/io_in_rdata_r[225] ;
wire \asic/lsdram/msdram/io_in_rdata_r[224] ;
wire \asic/lsdram/msdram/io_in_rdata_r[223] ;
wire \asic/lsdram/msdram/io_in_rdata_r[222] ;
wire \asic/lsdram/msdram/io_in_rdata_r[221] ;
wire \asic/lsdram/msdram/io_in_rdata_r[220] ;
wire \asic/lsdram/msdram/io_in_rdata_r[219] ;
wire \asic/lsdram/msdram/io_in_rdata_r[218] ;
wire \asic/lsdram/msdram/io_in_rdata_r[217] ;
wire \asic/lsdram/msdram/io_in_rdata_r[216] ;
wire \asic/lsdram/msdram/io_in_rdata_r[215] ;
wire \asic/lsdram/msdram/io_in_rdata_r[214] ;
wire \asic/lsdram/msdram/io_in_rdata_r[213] ;
wire \asic/lsdram/msdram/io_in_rdata_r[212] ;
wire \asic/lsdram/msdram/io_in_rdata_r[211] ;
wire \asic/lsdram/msdram/io_in_rdata_r[210] ;
wire \asic/lsdram/msdram/io_in_rdata_r[209] ;
wire \asic/lsdram/msdram/io_in_rdata_r[208] ;
wire \asic/lsdram/msdram/io_in_rdata_r[207] ;
wire \asic/lsdram/msdram/io_in_rdata_r[206] ;
wire \asic/lsdram/msdram/io_in_rdata_r[205] ;
wire \asic/lsdram/msdram/io_in_rdata_r[204] ;
wire \asic/lsdram/msdram/io_in_rdata_r[203] ;
wire \asic/lsdram/msdram/io_in_rdata_r[202] ;
wire \asic/lsdram/msdram/io_in_rdata_r[201] ;
wire \asic/lsdram/msdram/io_in_rdata_r[200] ;
wire \asic/lsdram/msdram/io_in_rdata_r[199] ;
wire \asic/lsdram/msdram/io_in_rdata_r[198] ;
wire \asic/lsdram/msdram/io_in_rdata_r[197] ;
wire \asic/lsdram/msdram/io_in_rdata_r[196] ;
wire \asic/lsdram/msdram/io_in_rdata_r[195] ;
wire \asic/lsdram/msdram/io_in_rdata_r[194] ;
wire \asic/lsdram/msdram/io_in_rdata_r[193] ;
wire \asic/lsdram/msdram/io_in_rdata_r[192] ;
wire \asic/lsdram/msdram/io_in_rdata_r[191] ;
wire \asic/lsdram/msdram/io_in_rdata_r[190] ;
wire \asic/lsdram/msdram/io_in_rdata_r[189] ;
wire \asic/lsdram/msdram/io_in_rdata_r[188] ;
wire \asic/lsdram/msdram/io_in_rdata_r[187] ;
wire \asic/lsdram/msdram/io_in_rdata_r[186] ;
wire \asic/lsdram/msdram/io_in_rdata_r[185] ;
wire \asic/lsdram/msdram/io_in_rdata_r[184] ;
wire \asic/lsdram/msdram/io_in_rdata_r[183] ;
wire \asic/lsdram/msdram/io_in_rdata_r[182] ;
wire \asic/lsdram/msdram/io_in_rdata_r[181] ;
wire \asic/lsdram/msdram/io_in_rdata_r[180] ;
wire \asic/lsdram/msdram/io_in_rdata_r[179] ;
wire \asic/lsdram/msdram/io_in_rdata_r[178] ;
wire \asic/lsdram/msdram/io_in_rdata_r[177] ;
wire \asic/lsdram/msdram/io_in_rdata_r[176] ;
wire \asic/lsdram/msdram/io_in_rdata_r[175] ;
wire \asic/lsdram/msdram/io_in_rdata_r[174] ;
wire \asic/lsdram/msdram/io_in_rdata_r[173] ;
wire \asic/lsdram/msdram/io_in_rdata_r[172] ;
wire \asic/lsdram/msdram/io_in_rdata_r[171] ;
wire \asic/lsdram/msdram/io_in_rdata_r[170] ;
wire \asic/lsdram/msdram/io_in_rdata_r[169] ;
wire \asic/lsdram/msdram/io_in_rdata_r[168] ;
wire \asic/lsdram/msdram/io_in_rdata_r[167] ;
wire \asic/lsdram/msdram/io_in_rdata_r[166] ;
wire \asic/lsdram/msdram/io_in_rdata_r[165] ;
wire \asic/lsdram/msdram/io_in_rdata_r[164] ;
wire \asic/lsdram/msdram/io_in_rdata_r[163] ;
wire \asic/lsdram/msdram/io_in_rdata_r[162] ;
wire \asic/lsdram/msdram/io_in_rdata_r[161] ;
wire \asic/lsdram/msdram/io_in_rdata_r[160] ;
wire \asic/lsdram/msdram/io_in_rdata_r[159] ;
wire \asic/lsdram/msdram/io_in_rdata_r[158] ;
wire \asic/lsdram/msdram/io_in_rdata_r[157] ;
wire \asic/lsdram/msdram/io_in_rdata_r[156] ;
wire \asic/lsdram/msdram/io_in_rdata_r[155] ;
wire \asic/lsdram/msdram/io_in_rdata_r[154] ;
wire \asic/lsdram/msdram/io_in_rdata_r[153] ;
wire \asic/lsdram/msdram/io_in_rdata_r[152] ;
wire \asic/lsdram/msdram/io_in_rdata_r[151] ;
wire \asic/lsdram/msdram/io_in_rdata_r[150] ;
wire \asic/lsdram/msdram/io_in_rdata_r[149] ;
wire \asic/lsdram/msdram/io_in_rdata_r[148] ;
wire \asic/lsdram/msdram/io_in_rdata_r[147] ;
wire \asic/lsdram/msdram/io_in_rdata_r[146] ;
wire \asic/lsdram/msdram/io_in_rdata_r[145] ;
wire \asic/lsdram/msdram/io_in_rdata_r[144] ;
wire \asic/lsdram/msdram/io_in_rdata_r[143] ;
wire \asic/lsdram/msdram/io_in_rdata_r[142] ;
wire \asic/lsdram/msdram/io_in_rdata_r[141] ;
wire \asic/lsdram/msdram/io_in_rdata_r[140] ;
wire \asic/lsdram/msdram/io_in_rdata_r[139] ;
wire \asic/lsdram/msdram/io_in_rdata_r[138] ;
wire \asic/lsdram/msdram/io_in_rdata_r[137] ;
wire \asic/lsdram/msdram/io_in_rdata_r[136] ;
wire \asic/lsdram/msdram/io_in_rdata_r[135] ;
wire \asic/lsdram/msdram/io_in_rdata_r[134] ;
wire \asic/lsdram/msdram/io_in_rdata_r[133] ;
wire \asic/lsdram/msdram/io_in_rdata_r[132] ;
wire \asic/lsdram/msdram/io_in_rdata_r[131] ;
wire \asic/lsdram/msdram/io_in_rdata_r[130] ;
wire \asic/lsdram/msdram/io_in_rdata_r[129] ;
wire \asic/lsdram/msdram/io_in_rdata_r[128] ;
wire \asic/lsdram/msdram/io_in_rdata_r[127] ;
wire \asic/lsdram/msdram/io_in_rdata_r[126] ;
wire \asic/lsdram/msdram/io_in_rdata_r[125] ;
wire \asic/lsdram/msdram/io_in_rdata_r[124] ;
wire \asic/lsdram/msdram/io_in_rdata_r[123] ;
wire \asic/lsdram/msdram/io_in_rdata_r[122] ;
wire \asic/lsdram/msdram/io_in_rdata_r[121] ;
wire \asic/lsdram/msdram/io_in_rdata_r[120] ;
wire \asic/lsdram/msdram/io_in_rdata_r[119] ;
wire \asic/lsdram/msdram/io_in_rdata_r[118] ;
wire \asic/lsdram/msdram/io_in_rdata_r[117] ;
wire \asic/lsdram/msdram/io_in_rdata_r[116] ;
wire \asic/lsdram/msdram/io_in_rdata_r[115] ;
wire \asic/lsdram/msdram/io_in_rdata_r[114] ;
wire \asic/lsdram/msdram/io_in_rdata_r[113] ;
wire \asic/lsdram/msdram/io_in_rdata_r[112] ;
wire \asic/lsdram/msdram/io_in_rdata_r[111] ;
wire \asic/lsdram/msdram/io_in_rdata_r[110] ;
wire \asic/lsdram/msdram/io_in_rdata_r[109] ;
wire \asic/lsdram/msdram/io_in_rdata_r[108] ;
wire \asic/lsdram/msdram/io_in_rdata_r[107] ;
wire \asic/lsdram/msdram/io_in_rdata_r[106] ;
wire \asic/lsdram/msdram/io_in_rdata_r[105] ;
wire \asic/lsdram/msdram/io_in_rdata_r[104] ;
wire \asic/lsdram/msdram/io_in_rdata_r[103] ;
wire \asic/lsdram/msdram/io_in_rdata_r[102] ;
wire \asic/lsdram/msdram/io_in_rdata_r[101] ;
wire \asic/lsdram/msdram/io_in_rdata_r[100] ;
wire \asic/lsdram/msdram/io_in_rdata_r[99] ;
wire \asic/lsdram/msdram/io_in_rdata_r[98] ;
wire \asic/lsdram/msdram/io_in_rdata_r[97] ;
wire \asic/lsdram/msdram/io_in_rdata_r[96] ;
wire \asic/lsdram/msdram/io_in_rdata_r[95] ;
wire \asic/lsdram/msdram/io_in_rdata_r[94] ;
wire \asic/lsdram/msdram/io_in_rdata_r[93] ;
wire \asic/lsdram/msdram/io_in_rdata_r[92] ;
wire \asic/lsdram/msdram/io_in_rdata_r[91] ;
wire \asic/lsdram/msdram/io_in_rdata_r[90] ;
wire \asic/lsdram/msdram/io_in_rdata_r[89] ;
wire \asic/lsdram/msdram/io_in_rdata_r[88] ;
wire \asic/lsdram/msdram/io_in_rdata_r[87] ;
wire \asic/lsdram/msdram/io_in_rdata_r[86] ;
wire \asic/lsdram/msdram/io_in_rdata_r[85] ;
wire \asic/lsdram/msdram/io_in_rdata_r[84] ;
wire \asic/lsdram/msdram/io_in_rdata_r[83] ;
wire \asic/lsdram/msdram/io_in_rdata_r[82] ;
wire \asic/lsdram/msdram/io_in_rdata_r[81] ;
wire \asic/lsdram/msdram/io_in_rdata_r[80] ;
wire \asic/lsdram/msdram/io_in_rdata_r[79] ;
wire \asic/lsdram/msdram/io_in_rdata_r[78] ;
wire \asic/lsdram/msdram/io_in_rdata_r[77] ;
wire \asic/lsdram/msdram/io_in_rdata_r[76] ;
wire \asic/lsdram/msdram/io_in_rdata_r[75] ;
wire \asic/lsdram/msdram/io_in_rdata_r[74] ;
wire \asic/lsdram/msdram/io_in_rdata_r[73] ;
wire \asic/lsdram/msdram/io_in_rdata_r[72] ;
wire \asic/lsdram/msdram/io_in_rdata_r[71] ;
wire \asic/lsdram/msdram/io_in_rdata_r[70] ;
wire \asic/lsdram/msdram/io_in_rdata_r[69] ;
wire \asic/lsdram/msdram/io_in_rdata_r[68] ;
wire \asic/lsdram/msdram/io_in_rdata_r[67] ;
wire \asic/lsdram/msdram/io_in_rdata_r[66] ;
wire \asic/lsdram/msdram/io_in_rdata_r[65] ;
wire \asic/lsdram/msdram/io_in_rdata_r[64] ;
wire \asic/lsdram/msdram/io_in_rdata_r[63] ;
wire \asic/lsdram/msdram/io_in_rdata_r[62] ;
wire \asic/lsdram/msdram/io_in_rdata_r[61] ;
wire \asic/lsdram/msdram/io_in_rdata_r[60] ;
wire \asic/lsdram/msdram/io_in_rdata_r[59] ;
wire \asic/lsdram/msdram/io_in_rdata_r[58] ;
wire \asic/lsdram/msdram/io_in_rdata_r[57] ;
wire \asic/lsdram/msdram/io_in_rdata_r[56] ;
wire \asic/lsdram/msdram/io_in_rdata_r[55] ;
wire \asic/lsdram/msdram/io_in_rdata_r[54] ;
wire \asic/lsdram/msdram/io_in_rdata_r[53] ;
wire \asic/lsdram/msdram/io_in_rdata_r[52] ;
wire \asic/lsdram/msdram/io_in_rdata_r[51] ;
wire \asic/lsdram/msdram/io_in_rdata_r[50] ;
wire \asic/lsdram/msdram/io_in_rdata_r[49] ;
wire \asic/lsdram/msdram/io_in_rdata_r[48] ;
wire \asic/lsdram/msdram/io_in_rdata_r[47] ;
wire \asic/lsdram/msdram/io_in_rdata_r[46] ;
wire \asic/lsdram/msdram/io_in_rdata_r[45] ;
wire \asic/lsdram/msdram/io_in_rdata_r[44] ;
wire \asic/lsdram/msdram/io_in_rdata_r[43] ;
wire \asic/lsdram/msdram/io_in_rdata_r[42] ;
wire \asic/lsdram/msdram/io_in_rdata_r[41] ;
wire \asic/lsdram/msdram/io_in_rdata_r[40] ;
wire \asic/lsdram/msdram/io_in_rdata_r[39] ;
wire \asic/lsdram/msdram/io_in_rdata_r[38] ;
wire \asic/lsdram/msdram/io_in_rdata_r[37] ;
wire \asic/lsdram/msdram/io_in_rdata_r[36] ;
wire \asic/lsdram/msdram/io_in_rdata_r[35] ;
wire \asic/lsdram/msdram/io_in_rdata_r[34] ;
wire \asic/lsdram/msdram/io_in_rdata_r[33] ;
wire \asic/lsdram/msdram/io_in_rdata_r[32] ;
wire \asic/lsdram/msdram/io_in_rdata_r[31] ;
wire \asic/lsdram/msdram/io_in_rdata_r[30] ;
wire \asic/lsdram/msdram/io_in_rdata_r[29] ;
wire \asic/lsdram/msdram/io_in_rdata_r[28] ;
wire \asic/lsdram/msdram/io_in_rdata_r[27] ;
wire \asic/lsdram/msdram/io_in_rdata_r[26] ;
wire \asic/lsdram/msdram/io_in_rdata_r[25] ;
wire \asic/lsdram/msdram/io_in_rdata_r[24] ;
wire \asic/lsdram/msdram/io_in_rdata_r[23] ;
wire \asic/lsdram/msdram/io_in_rdata_r[22] ;
wire \asic/lsdram/msdram/io_in_rdata_r[21] ;
wire \asic/lsdram/msdram/io_in_rdata_r[20] ;
wire \asic/lsdram/msdram/io_in_rdata_r[19] ;
wire \asic/lsdram/msdram/io_in_rdata_r[18] ;
wire \asic/lsdram/msdram/io_in_rdata_r[17] ;
wire \asic/lsdram/msdram/io_in_rdata_r[16] ;
wire \asic/lsdram/msdram/io_in_rdata_r[15] ;
wire \asic/lsdram/msdram/io_in_rdata_r[14] ;
wire \asic/lsdram/msdram/io_in_rdata_r[13] ;
wire \asic/lsdram/msdram/io_in_rdata_r[12] ;
wire \asic/lsdram/msdram/io_in_rdata_r[11] ;
wire \asic/lsdram/msdram/io_in_rdata_r[10] ;
wire \asic/lsdram/msdram/io_in_rdata_r[9] ;
wire \asic/lsdram/msdram/io_in_rdata_r[8] ;
wire \asic/lsdram/msdram/io_in_rdata_r[7] ;
wire \asic/lsdram/msdram/io_in_rdata_r[6] ;
wire \asic/lsdram/msdram/io_in_rdata_r[5] ;
wire \asic/lsdram/msdram/io_in_rdata_r[4] ;
wire \asic/lsdram/msdram/io_in_rdata_r[3] ;
wire \asic/lsdram/msdram/io_in_rdata_r[2] ;
wire \asic/lsdram/msdram/io_in_rdata_r[1] ;
wire \asic/lsdram/msdram/io_in_rdata_r[0] ;
wire \asic/lsdram/msdram/io_clk_out ;
wire \asic/lsdram/msdram/io_in_awready ;
wire \asic/lsdram/msdram/io_in_awvalid ;
wire \asic/lsdram/msdram/io_in_wready ;
wire \asic/lsdram/msdram/io_in_wvalid ;
wire \asic/lsdram/msdram/io_in_bready ;
wire \asic/lsdram/msdram/io_in_bvalid ;
wire \asic/lsdram/msdram/io_in_arready ;
wire \asic/lsdram/msdram/io_in_arvalid ;
wire \asic/lsdram/msdram/io_in_rready ;
wire \asic/lsdram/msdram/io_in_rvalid ;
wire \asic/lsdram/msdram/io_dmi_cmd_en ;
wire \asic/lsdram/msdram/io_dmi_wr_data_en ;
wire \asic/lsdram/msdram/io_dmi_wr_data_end ;
wire \asic/lsdram/msdram/io_dmi_clk_out ;
wire \asic/lsdram/msdram/io_dmi_init_calib_complete ;
wire \asic/lsdram/msdram/io_dmi_cmd_ready ;
wire \asic/lsdram/msdram/io_dmi_wr_data_rdy ;
wire \asic/lsdram/msdram/io_dmi_rd_data_valid ;
wire clock;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\asic/cpu/cpu/if_stage/fs_pc[31] ,\asic/cpu/cpu/if_stage/fs_pc[30] ,\asic/cpu/cpu/if_stage/fs_pc[29] ,\asic/cpu/cpu/if_stage/fs_pc[28] ,\asic/cpu/cpu/if_stage/fs_pc[27] ,\asic/cpu/cpu/if_stage/fs_pc[26] ,\asic/cpu/cpu/if_stage/fs_pc[25] ,\asic/cpu/cpu/if_stage/fs_pc[24] ,\asic/cpu/cpu/if_stage/fs_pc[23] ,\asic/cpu/cpu/if_stage/fs_pc[22] ,\asic/cpu/cpu/if_stage/fs_pc[21] ,\asic/cpu/cpu/if_stage/fs_pc[20] ,\asic/cpu/cpu/if_stage/fs_pc[19] ,\asic/cpu/cpu/if_stage/fs_pc[18] ,\asic/cpu/cpu/if_stage/fs_pc[17] ,\asic/cpu/cpu/if_stage/fs_pc[16] ,\asic/cpu/cpu/if_stage/fs_pc[15] ,\asic/cpu/cpu/if_stage/fs_pc[14] ,\asic/cpu/cpu/if_stage/fs_pc[13] ,\asic/cpu/cpu/if_stage/fs_pc[12] ,\asic/cpu/cpu/if_stage/fs_pc[11] ,\asic/cpu/cpu/if_stage/fs_pc[10] ,\asic/cpu/cpu/if_stage/fs_pc[9] ,\asic/cpu/cpu/if_stage/fs_pc[8] ,\asic/cpu/cpu/if_stage/fs_pc[7] ,\asic/cpu/cpu/if_stage/fs_pc[6] ,\asic/cpu/cpu/if_stage/fs_pc[5] ,\asic/cpu/cpu/if_stage/fs_pc[4] ,\asic/cpu/cpu/if_stage/fs_pc[3] ,\asic/cpu/cpu/if_stage/fs_pc[2] ,\asic/cpu/cpu/if_stage/fs_pc[1] ,\asic/cpu/cpu/if_stage/fs_pc[0] }),
    .data_i({\asic/cpu/cpu/if_stage/fs_pc[31] ,\asic/cpu/cpu/if_stage/fs_pc[30] ,\asic/cpu/cpu/if_stage/fs_pc[29] ,\asic/cpu/cpu/if_stage/fs_pc[28] ,\asic/cpu/cpu/if_stage/fs_pc[27] ,\asic/cpu/cpu/if_stage/fs_pc[26] ,\asic/cpu/cpu/if_stage/fs_pc[25] ,\asic/cpu/cpu/if_stage/fs_pc[24] ,\asic/cpu/cpu/if_stage/fs_pc[23] ,\asic/cpu/cpu/if_stage/fs_pc[22] ,\asic/cpu/cpu/if_stage/fs_pc[21] ,\asic/cpu/cpu/if_stage/fs_pc[20] ,\asic/cpu/cpu/if_stage/fs_pc[19] ,\asic/cpu/cpu/if_stage/fs_pc[18] ,\asic/cpu/cpu/if_stage/fs_pc[17] ,\asic/cpu/cpu/if_stage/fs_pc[16] ,\asic/cpu/cpu/if_stage/fs_pc[15] ,\asic/cpu/cpu/if_stage/fs_pc[14] ,\asic/cpu/cpu/if_stage/fs_pc[13] ,\asic/cpu/cpu/if_stage/fs_pc[12] ,\asic/cpu/cpu/if_stage/fs_pc[11] ,\asic/cpu/cpu/if_stage/fs_pc[10] ,\asic/cpu/cpu/if_stage/fs_pc[9] ,\asic/cpu/cpu/if_stage/fs_pc[8] ,\asic/cpu/cpu/if_stage/fs_pc[7] ,\asic/cpu/cpu/if_stage/fs_pc[6] ,\asic/cpu/cpu/if_stage/fs_pc[5] ,\asic/cpu/cpu/if_stage/fs_pc[4] ,\asic/cpu/cpu/if_stage/fs_pc[3] ,\asic/cpu/cpu/if_stage/fs_pc[2] ,\asic/cpu/cpu/if_stage/fs_pc[1] ,\asic/cpu/cpu/if_stage/fs_pc[0] ,\asic/cpu/cpu/if_stage/fs_inst[31] ,\asic/cpu/cpu/if_stage/fs_inst[30] ,\asic/cpu/cpu/if_stage/fs_inst[29] ,\asic/cpu/cpu/if_stage/fs_inst[28] ,\asic/cpu/cpu/if_stage/fs_inst[27] ,\asic/cpu/cpu/if_stage/fs_inst[26] ,\asic/cpu/cpu/if_stage/fs_inst[25] ,\asic/cpu/cpu/if_stage/fs_inst[24] ,\asic/cpu/cpu/if_stage/fs_inst[23] ,\asic/cpu/cpu/if_stage/fs_inst[22] ,\asic/cpu/cpu/if_stage/fs_inst[21] ,\asic/cpu/cpu/if_stage/fs_inst[20] ,\asic/cpu/cpu/if_stage/fs_inst[19] ,\asic/cpu/cpu/if_stage/fs_inst[18] ,\asic/cpu/cpu/if_stage/fs_inst[17] ,\asic/cpu/cpu/if_stage/fs_inst[16] ,\asic/cpu/cpu/if_stage/fs_inst[15] ,\asic/cpu/cpu/if_stage/fs_inst[14] ,\asic/cpu/cpu/if_stage/fs_inst[13] ,\asic/cpu/cpu/if_stage/fs_inst[12] ,\asic/cpu/cpu/if_stage/fs_inst[11] ,\asic/cpu/cpu/if_stage/fs_inst[10] ,\asic/cpu/cpu/if_stage/fs_inst[9] ,\asic/cpu/cpu/if_stage/fs_inst[8] ,\asic/cpu/cpu/if_stage/fs_inst[7] ,\asic/cpu/cpu/if_stage/fs_inst[6] ,\asic/cpu/cpu/if_stage/fs_inst[5] ,\asic/cpu/cpu/if_stage/fs_inst[4] ,\asic/cpu/cpu/if_stage/fs_inst[3] ,\asic/cpu/cpu/if_stage/fs_inst[2] ,\asic/cpu/cpu/if_stage/fs_inst[1] ,\asic/cpu/cpu/if_stage/fs_inst[0] ,\asic/lsdram/msdram/io_in_awid[3] ,\asic/lsdram/msdram/io_in_awid[2] ,\asic/lsdram/msdram/io_in_awid[1] ,\asic/lsdram/msdram/io_in_awid[0] ,\asic/lsdram/msdram/io_in_awaddr[31] ,\asic/lsdram/msdram/io_in_awaddr[30] ,\asic/lsdram/msdram/io_in_awaddr[29] ,\asic/lsdram/msdram/io_in_awaddr[28] ,\asic/lsdram/msdram/io_in_awaddr[27] ,\asic/lsdram/msdram/io_in_awaddr[26] ,\asic/lsdram/msdram/io_in_awaddr[25] ,\asic/lsdram/msdram/io_in_awaddr[24] ,\asic/lsdram/msdram/io_in_awaddr[23] ,\asic/lsdram/msdram/io_in_awaddr[22] ,\asic/lsdram/msdram/io_in_awaddr[21] ,\asic/lsdram/msdram/io_in_awaddr[20] ,\asic/lsdram/msdram/io_in_awaddr[19] ,\asic/lsdram/msdram/io_in_awaddr[18] ,\asic/lsdram/msdram/io_in_awaddr[17] ,\asic/lsdram/msdram/io_in_awaddr[16] ,\asic/lsdram/msdram/io_in_awaddr[15] ,\asic/lsdram/msdram/io_in_awaddr[14] ,\asic/lsdram/msdram/io_in_awaddr[13] ,\asic/lsdram/msdram/io_in_awaddr[12] ,\asic/lsdram/msdram/io_in_awaddr[11] ,\asic/lsdram/msdram/io_in_awaddr[10] ,\asic/lsdram/msdram/io_in_awaddr[9] ,\asic/lsdram/msdram/io_in_awaddr[8] ,\asic/lsdram/msdram/io_in_awaddr[7] ,\asic/lsdram/msdram/io_in_awaddr[6] ,\asic/lsdram/msdram/io_in_awaddr[5] ,\asic/lsdram/msdram/io_in_awaddr[4] ,\asic/lsdram/msdram/io_in_awaddr[3] ,\asic/lsdram/msdram/io_in_awaddr[2] ,\asic/lsdram/msdram/io_in_awaddr[1] ,\asic/lsdram/msdram/io_in_awaddr[0] ,\asic/lsdram/msdram/io_in_awlen[7] ,\asic/lsdram/msdram/io_in_awlen[6] ,\asic/lsdram/msdram/io_in_awlen[5] ,\asic/lsdram/msdram/io_in_awlen[4] ,\asic/lsdram/msdram/io_in_awlen[3] ,\asic/lsdram/msdram/io_in_awlen[2] ,\asic/lsdram/msdram/io_in_awlen[1] ,\asic/lsdram/msdram/io_in_awlen[0] ,\asic/lsdram/msdram/io_in_awsize[2] ,\asic/lsdram/msdram/io_in_awsize[1] ,\asic/lsdram/msdram/io_in_awsize[0] ,\asic/lsdram/msdram/io_in_wdata[31] ,\asic/lsdram/msdram/io_in_wdata[30] ,\asic/lsdram/msdram/io_in_wdata[29] ,\asic/lsdram/msdram/io_in_wdata[28] ,\asic/lsdram/msdram/io_in_wdata[27] ,\asic/lsdram/msdram/io_in_wdata[26] ,\asic/lsdram/msdram/io_in_wdata[25] ,\asic/lsdram/msdram/io_in_wdata[24] ,\asic/lsdram/msdram/io_in_wdata[23] ,\asic/lsdram/msdram/io_in_wdata[22] ,\asic/lsdram/msdram/io_in_wdata[21] ,\asic/lsdram/msdram/io_in_wdata[20] ,\asic/lsdram/msdram/io_in_wdata[19] ,\asic/lsdram/msdram/io_in_wdata[18] ,\asic/lsdram/msdram/io_in_wdata[17] ,\asic/lsdram/msdram/io_in_wdata[16] ,\asic/lsdram/msdram/io_in_wdata[15] ,\asic/lsdram/msdram/io_in_wdata[14] ,\asic/lsdram/msdram/io_in_wdata[13] ,\asic/lsdram/msdram/io_in_wdata[12] ,\asic/lsdram/msdram/io_in_wdata[11] ,\asic/lsdram/msdram/io_in_wdata[10] ,\asic/lsdram/msdram/io_in_wdata[9] ,\asic/lsdram/msdram/io_in_wdata[8] ,\asic/lsdram/msdram/io_in_wdata[7] ,\asic/lsdram/msdram/io_in_wdata[6] ,\asic/lsdram/msdram/io_in_wdata[5] ,\asic/lsdram/msdram/io_in_wdata[4] ,\asic/lsdram/msdram/io_in_wdata[3] ,\asic/lsdram/msdram/io_in_wdata[2] ,\asic/lsdram/msdram/io_in_wdata[1] ,\asic/lsdram/msdram/io_in_wdata[0] ,\asic/lsdram/msdram/io_in_wstrb[3] ,\asic/lsdram/msdram/io_in_wstrb[2] ,\asic/lsdram/msdram/io_in_wstrb[1] ,\asic/lsdram/msdram/io_in_wstrb[0] ,\asic/lsdram/msdram/io_in_bid[3] ,\asic/lsdram/msdram/io_in_bid[2] ,\asic/lsdram/msdram/io_in_bid[1] ,\asic/lsdram/msdram/io_in_bid[0] ,\asic/lsdram/msdram/io_in_arid[3] ,\asic/lsdram/msdram/io_in_arid[2] ,\asic/lsdram/msdram/io_in_arid[1] ,\asic/lsdram/msdram/io_in_arid[0] ,\asic/lsdram/msdram/io_in_araddr[31] ,\asic/lsdram/msdram/io_in_araddr[30] ,\asic/lsdram/msdram/io_in_araddr[29] ,\asic/lsdram/msdram/io_in_araddr[28] ,\asic/lsdram/msdram/io_in_araddr[27] ,\asic/lsdram/msdram/io_in_araddr[26] ,\asic/lsdram/msdram/io_in_araddr[25] ,\asic/lsdram/msdram/io_in_araddr[24] ,\asic/lsdram/msdram/io_in_araddr[23] ,\asic/lsdram/msdram/io_in_araddr[22] ,\asic/lsdram/msdram/io_in_araddr[21] ,\asic/lsdram/msdram/io_in_araddr[20] ,\asic/lsdram/msdram/io_in_araddr[19] ,\asic/lsdram/msdram/io_in_araddr[18] ,\asic/lsdram/msdram/io_in_araddr[17] ,\asic/lsdram/msdram/io_in_araddr[16] ,\asic/lsdram/msdram/io_in_araddr[15] ,\asic/lsdram/msdram/io_in_araddr[14] ,\asic/lsdram/msdram/io_in_araddr[13] ,\asic/lsdram/msdram/io_in_araddr[12] ,\asic/lsdram/msdram/io_in_araddr[11] ,\asic/lsdram/msdram/io_in_araddr[10] ,\asic/lsdram/msdram/io_in_araddr[9] ,\asic/lsdram/msdram/io_in_araddr[8] ,\asic/lsdram/msdram/io_in_araddr[7] ,\asic/lsdram/msdram/io_in_araddr[6] ,\asic/lsdram/msdram/io_in_araddr[5] ,\asic/lsdram/msdram/io_in_araddr[4] ,\asic/lsdram/msdram/io_in_araddr[3] ,\asic/lsdram/msdram/io_in_araddr[2] ,\asic/lsdram/msdram/io_in_araddr[1] ,\asic/lsdram/msdram/io_in_araddr[0] ,\asic/lsdram/msdram/io_in_arlen[7] ,\asic/lsdram/msdram/io_in_arlen[6] ,\asic/lsdram/msdram/io_in_arlen[5] ,\asic/lsdram/msdram/io_in_arlen[4] ,\asic/lsdram/msdram/io_in_arlen[3] ,\asic/lsdram/msdram/io_in_arlen[2] ,\asic/lsdram/msdram/io_in_arlen[1] ,\asic/lsdram/msdram/io_in_arlen[0] ,\asic/lsdram/msdram/io_in_arsize[2] ,\asic/lsdram/msdram/io_in_arsize[1] ,\asic/lsdram/msdram/io_in_arsize[0] ,\asic/lsdram/msdram/io_in_rid[3] ,\asic/lsdram/msdram/io_in_rid[2] ,\asic/lsdram/msdram/io_in_rid[1] ,\asic/lsdram/msdram/io_in_rid[0] ,\asic/lsdram/msdram/io_in_rdata[31] ,\asic/lsdram/msdram/io_in_rdata[30] ,\asic/lsdram/msdram/io_in_rdata[29] ,\asic/lsdram/msdram/io_in_rdata[28] ,\asic/lsdram/msdram/io_in_rdata[27] ,\asic/lsdram/msdram/io_in_rdata[26] ,\asic/lsdram/msdram/io_in_rdata[25] ,\asic/lsdram/msdram/io_in_rdata[24] ,\asic/lsdram/msdram/io_in_rdata[23] ,\asic/lsdram/msdram/io_in_rdata[22] ,\asic/lsdram/msdram/io_in_rdata[21] ,\asic/lsdram/msdram/io_in_rdata[20] ,\asic/lsdram/msdram/io_in_rdata[19] ,\asic/lsdram/msdram/io_in_rdata[18] ,\asic/lsdram/msdram/io_in_rdata[17] ,\asic/lsdram/msdram/io_in_rdata[16] ,\asic/lsdram/msdram/io_in_rdata[15] ,\asic/lsdram/msdram/io_in_rdata[14] ,\asic/lsdram/msdram/io_in_rdata[13] ,\asic/lsdram/msdram/io_in_rdata[12] ,\asic/lsdram/msdram/io_in_rdata[11] ,\asic/lsdram/msdram/io_in_rdata[10] ,\asic/lsdram/msdram/io_in_rdata[9] ,\asic/lsdram/msdram/io_in_rdata[8] ,\asic/lsdram/msdram/io_in_rdata[7] ,\asic/lsdram/msdram/io_in_rdata[6] ,\asic/lsdram/msdram/io_in_rdata[5] ,\asic/lsdram/msdram/io_in_rdata[4] ,\asic/lsdram/msdram/io_in_rdata[3] ,\asic/lsdram/msdram/io_in_rdata[2] ,\asic/lsdram/msdram/io_in_rdata[1] ,\asic/lsdram/msdram/io_in_rdata[0] ,\asic/lsdram/msdram/io_dmi_cmd[2] ,\asic/lsdram/msdram/io_dmi_cmd[1] ,\asic/lsdram/msdram/io_dmi_cmd[0] ,\asic/lsdram/msdram/io_dmi_addr[28] ,\asic/lsdram/msdram/io_dmi_addr[27] ,\asic/lsdram/msdram/io_dmi_addr[26] ,\asic/lsdram/msdram/io_dmi_addr[25] ,\asic/lsdram/msdram/io_dmi_addr[24] ,\asic/lsdram/msdram/io_dmi_addr[23] ,\asic/lsdram/msdram/io_dmi_addr[22] ,\asic/lsdram/msdram/io_dmi_addr[21] ,\asic/lsdram/msdram/io_dmi_addr[20] ,\asic/lsdram/msdram/io_dmi_addr[19] ,\asic/lsdram/msdram/io_dmi_addr[18] ,\asic/lsdram/msdram/io_dmi_addr[17] ,\asic/lsdram/msdram/io_dmi_addr[16] ,\asic/lsdram/msdram/io_dmi_addr[15] ,\asic/lsdram/msdram/io_dmi_addr[14] ,\asic/lsdram/msdram/io_dmi_addr[13] ,\asic/lsdram/msdram/io_dmi_addr[12] ,\asic/lsdram/msdram/io_dmi_addr[11] ,\asic/lsdram/msdram/io_dmi_addr[10] ,\asic/lsdram/msdram/io_dmi_addr[9] ,\asic/lsdram/msdram/io_dmi_addr[8] ,\asic/lsdram/msdram/io_dmi_addr[7] ,\asic/lsdram/msdram/io_dmi_addr[6] ,\asic/lsdram/msdram/io_dmi_addr[5] ,\asic/lsdram/msdram/io_dmi_addr[4] ,\asic/lsdram/msdram/io_dmi_addr[3] ,\asic/lsdram/msdram/io_dmi_addr[2] ,\asic/lsdram/msdram/io_dmi_addr[1] ,\asic/lsdram/msdram/io_dmi_addr[0] ,\asic/lsdram/msdram/io_dmi_wr_data[255] ,\asic/lsdram/msdram/io_dmi_wr_data[254] ,\asic/lsdram/msdram/io_dmi_wr_data[253] ,\asic/lsdram/msdram/io_dmi_wr_data[252] ,\asic/lsdram/msdram/io_dmi_wr_data[251] ,\asic/lsdram/msdram/io_dmi_wr_data[250] ,\asic/lsdram/msdram/io_dmi_wr_data[249] ,\asic/lsdram/msdram/io_dmi_wr_data[248] ,\asic/lsdram/msdram/io_dmi_wr_data[247] ,\asic/lsdram/msdram/io_dmi_wr_data[246] ,\asic/lsdram/msdram/io_dmi_wr_data[245] ,\asic/lsdram/msdram/io_dmi_wr_data[244] ,\asic/lsdram/msdram/io_dmi_wr_data[243] ,\asic/lsdram/msdram/io_dmi_wr_data[242] ,\asic/lsdram/msdram/io_dmi_wr_data[241] ,\asic/lsdram/msdram/io_dmi_wr_data[240] ,\asic/lsdram/msdram/io_dmi_wr_data[239] ,\asic/lsdram/msdram/io_dmi_wr_data[238] ,\asic/lsdram/msdram/io_dmi_wr_data[237] ,\asic/lsdram/msdram/io_dmi_wr_data[236] ,\asic/lsdram/msdram/io_dmi_wr_data[235] ,\asic/lsdram/msdram/io_dmi_wr_data[234] ,\asic/lsdram/msdram/io_dmi_wr_data[233] ,\asic/lsdram/msdram/io_dmi_wr_data[232] ,\asic/lsdram/msdram/io_dmi_wr_data[231] ,\asic/lsdram/msdram/io_dmi_wr_data[230] ,\asic/lsdram/msdram/io_dmi_wr_data[229] ,\asic/lsdram/msdram/io_dmi_wr_data[228] ,\asic/lsdram/msdram/io_dmi_wr_data[227] ,\asic/lsdram/msdram/io_dmi_wr_data[226] ,\asic/lsdram/msdram/io_dmi_wr_data[225] ,\asic/lsdram/msdram/io_dmi_wr_data[224] ,\asic/lsdram/msdram/io_dmi_wr_data[223] ,\asic/lsdram/msdram/io_dmi_wr_data[222] ,\asic/lsdram/msdram/io_dmi_wr_data[221] ,\asic/lsdram/msdram/io_dmi_wr_data[220] ,\asic/lsdram/msdram/io_dmi_wr_data[219] ,\asic/lsdram/msdram/io_dmi_wr_data[218] ,\asic/lsdram/msdram/io_dmi_wr_data[217] ,\asic/lsdram/msdram/io_dmi_wr_data[216] ,\asic/lsdram/msdram/io_dmi_wr_data[215] ,\asic/lsdram/msdram/io_dmi_wr_data[214] ,\asic/lsdram/msdram/io_dmi_wr_data[213] ,\asic/lsdram/msdram/io_dmi_wr_data[212] ,\asic/lsdram/msdram/io_dmi_wr_data[211] ,\asic/lsdram/msdram/io_dmi_wr_data[210] ,\asic/lsdram/msdram/io_dmi_wr_data[209] ,\asic/lsdram/msdram/io_dmi_wr_data[208] ,\asic/lsdram/msdram/io_dmi_wr_data[207] ,\asic/lsdram/msdram/io_dmi_wr_data[206] ,\asic/lsdram/msdram/io_dmi_wr_data[205] ,\asic/lsdram/msdram/io_dmi_wr_data[204] ,\asic/lsdram/msdram/io_dmi_wr_data[203] ,\asic/lsdram/msdram/io_dmi_wr_data[202] ,\asic/lsdram/msdram/io_dmi_wr_data[201] ,\asic/lsdram/msdram/io_dmi_wr_data[200] ,\asic/lsdram/msdram/io_dmi_wr_data[199] ,\asic/lsdram/msdram/io_dmi_wr_data[198] ,\asic/lsdram/msdram/io_dmi_wr_data[197] ,\asic/lsdram/msdram/io_dmi_wr_data[196] ,\asic/lsdram/msdram/io_dmi_wr_data[195] ,\asic/lsdram/msdram/io_dmi_wr_data[194] ,\asic/lsdram/msdram/io_dmi_wr_data[193] ,\asic/lsdram/msdram/io_dmi_wr_data[192] ,\asic/lsdram/msdram/io_dmi_wr_data[191] ,\asic/lsdram/msdram/io_dmi_wr_data[190] ,\asic/lsdram/msdram/io_dmi_wr_data[189] ,\asic/lsdram/msdram/io_dmi_wr_data[188] ,\asic/lsdram/msdram/io_dmi_wr_data[187] ,\asic/lsdram/msdram/io_dmi_wr_data[186] ,\asic/lsdram/msdram/io_dmi_wr_data[185] ,\asic/lsdram/msdram/io_dmi_wr_data[184] ,\asic/lsdram/msdram/io_dmi_wr_data[183] ,\asic/lsdram/msdram/io_dmi_wr_data[182] ,\asic/lsdram/msdram/io_dmi_wr_data[181] ,\asic/lsdram/msdram/io_dmi_wr_data[180] ,\asic/lsdram/msdram/io_dmi_wr_data[179] ,\asic/lsdram/msdram/io_dmi_wr_data[178] ,\asic/lsdram/msdram/io_dmi_wr_data[177] ,\asic/lsdram/msdram/io_dmi_wr_data[176] ,\asic/lsdram/msdram/io_dmi_wr_data[175] ,\asic/lsdram/msdram/io_dmi_wr_data[174] ,\asic/lsdram/msdram/io_dmi_wr_data[173] ,\asic/lsdram/msdram/io_dmi_wr_data[172] ,\asic/lsdram/msdram/io_dmi_wr_data[171] ,\asic/lsdram/msdram/io_dmi_wr_data[170] ,\asic/lsdram/msdram/io_dmi_wr_data[169] ,\asic/lsdram/msdram/io_dmi_wr_data[168] ,\asic/lsdram/msdram/io_dmi_wr_data[167] ,\asic/lsdram/msdram/io_dmi_wr_data[166] ,\asic/lsdram/msdram/io_dmi_wr_data[165] ,\asic/lsdram/msdram/io_dmi_wr_data[164] ,\asic/lsdram/msdram/io_dmi_wr_data[163] ,\asic/lsdram/msdram/io_dmi_wr_data[162] ,\asic/lsdram/msdram/io_dmi_wr_data[161] ,\asic/lsdram/msdram/io_dmi_wr_data[160] ,\asic/lsdram/msdram/io_dmi_wr_data[159] ,\asic/lsdram/msdram/io_dmi_wr_data[158] ,\asic/lsdram/msdram/io_dmi_wr_data[157] ,\asic/lsdram/msdram/io_dmi_wr_data[156] ,\asic/lsdram/msdram/io_dmi_wr_data[155] ,\asic/lsdram/msdram/io_dmi_wr_data[154] ,\asic/lsdram/msdram/io_dmi_wr_data[153] ,\asic/lsdram/msdram/io_dmi_wr_data[152] ,\asic/lsdram/msdram/io_dmi_wr_data[151] ,\asic/lsdram/msdram/io_dmi_wr_data[150] ,\asic/lsdram/msdram/io_dmi_wr_data[149] ,\asic/lsdram/msdram/io_dmi_wr_data[148] ,\asic/lsdram/msdram/io_dmi_wr_data[147] ,\asic/lsdram/msdram/io_dmi_wr_data[146] ,\asic/lsdram/msdram/io_dmi_wr_data[145] ,\asic/lsdram/msdram/io_dmi_wr_data[144] ,\asic/lsdram/msdram/io_dmi_wr_data[143] ,\asic/lsdram/msdram/io_dmi_wr_data[142] ,\asic/lsdram/msdram/io_dmi_wr_data[141] ,\asic/lsdram/msdram/io_dmi_wr_data[140] ,\asic/lsdram/msdram/io_dmi_wr_data[139] ,\asic/lsdram/msdram/io_dmi_wr_data[138] ,\asic/lsdram/msdram/io_dmi_wr_data[137] ,\asic/lsdram/msdram/io_dmi_wr_data[136] ,\asic/lsdram/msdram/io_dmi_wr_data[135] ,\asic/lsdram/msdram/io_dmi_wr_data[134] ,\asic/lsdram/msdram/io_dmi_wr_data[133] ,\asic/lsdram/msdram/io_dmi_wr_data[132] ,\asic/lsdram/msdram/io_dmi_wr_data[131] ,\asic/lsdram/msdram/io_dmi_wr_data[130] ,\asic/lsdram/msdram/io_dmi_wr_data[129] ,\asic/lsdram/msdram/io_dmi_wr_data[128] ,\asic/lsdram/msdram/io_dmi_wr_data[127] ,\asic/lsdram/msdram/io_dmi_wr_data[126] ,\asic/lsdram/msdram/io_dmi_wr_data[125] ,\asic/lsdram/msdram/io_dmi_wr_data[124] ,\asic/lsdram/msdram/io_dmi_wr_data[123] ,\asic/lsdram/msdram/io_dmi_wr_data[122] ,\asic/lsdram/msdram/io_dmi_wr_data[121] ,\asic/lsdram/msdram/io_dmi_wr_data[120] ,\asic/lsdram/msdram/io_dmi_wr_data[119] ,\asic/lsdram/msdram/io_dmi_wr_data[118] ,\asic/lsdram/msdram/io_dmi_wr_data[117] ,\asic/lsdram/msdram/io_dmi_wr_data[116] ,\asic/lsdram/msdram/io_dmi_wr_data[115] ,\asic/lsdram/msdram/io_dmi_wr_data[114] ,\asic/lsdram/msdram/io_dmi_wr_data[113] ,\asic/lsdram/msdram/io_dmi_wr_data[112] ,\asic/lsdram/msdram/io_dmi_wr_data[111] ,\asic/lsdram/msdram/io_dmi_wr_data[110] ,\asic/lsdram/msdram/io_dmi_wr_data[109] ,\asic/lsdram/msdram/io_dmi_wr_data[108] ,\asic/lsdram/msdram/io_dmi_wr_data[107] ,\asic/lsdram/msdram/io_dmi_wr_data[106] ,\asic/lsdram/msdram/io_dmi_wr_data[105] ,\asic/lsdram/msdram/io_dmi_wr_data[104] ,\asic/lsdram/msdram/io_dmi_wr_data[103] ,\asic/lsdram/msdram/io_dmi_wr_data[102] ,\asic/lsdram/msdram/io_dmi_wr_data[101] ,\asic/lsdram/msdram/io_dmi_wr_data[100] ,\asic/lsdram/msdram/io_dmi_wr_data[99] ,\asic/lsdram/msdram/io_dmi_wr_data[98] ,\asic/lsdram/msdram/io_dmi_wr_data[97] ,\asic/lsdram/msdram/io_dmi_wr_data[96] ,\asic/lsdram/msdram/io_dmi_wr_data[95] ,\asic/lsdram/msdram/io_dmi_wr_data[94] ,\asic/lsdram/msdram/io_dmi_wr_data[93] ,\asic/lsdram/msdram/io_dmi_wr_data[92] ,\asic/lsdram/msdram/io_dmi_wr_data[91] ,\asic/lsdram/msdram/io_dmi_wr_data[90] ,\asic/lsdram/msdram/io_dmi_wr_data[89] ,\asic/lsdram/msdram/io_dmi_wr_data[88] ,\asic/lsdram/msdram/io_dmi_wr_data[87] ,\asic/lsdram/msdram/io_dmi_wr_data[86] ,\asic/lsdram/msdram/io_dmi_wr_data[85] ,\asic/lsdram/msdram/io_dmi_wr_data[84] ,\asic/lsdram/msdram/io_dmi_wr_data[83] ,\asic/lsdram/msdram/io_dmi_wr_data[82] ,\asic/lsdram/msdram/io_dmi_wr_data[81] ,\asic/lsdram/msdram/io_dmi_wr_data[80] ,\asic/lsdram/msdram/io_dmi_wr_data[79] ,\asic/lsdram/msdram/io_dmi_wr_data[78] ,\asic/lsdram/msdram/io_dmi_wr_data[77] ,\asic/lsdram/msdram/io_dmi_wr_data[76] ,\asic/lsdram/msdram/io_dmi_wr_data[75] ,\asic/lsdram/msdram/io_dmi_wr_data[74] ,\asic/lsdram/msdram/io_dmi_wr_data[73] ,\asic/lsdram/msdram/io_dmi_wr_data[72] ,\asic/lsdram/msdram/io_dmi_wr_data[71] ,\asic/lsdram/msdram/io_dmi_wr_data[70] ,\asic/lsdram/msdram/io_dmi_wr_data[69] ,\asic/lsdram/msdram/io_dmi_wr_data[68] ,\asic/lsdram/msdram/io_dmi_wr_data[67] ,\asic/lsdram/msdram/io_dmi_wr_data[66] ,\asic/lsdram/msdram/io_dmi_wr_data[65] ,\asic/lsdram/msdram/io_dmi_wr_data[64] ,\asic/lsdram/msdram/io_dmi_wr_data[63] ,\asic/lsdram/msdram/io_dmi_wr_data[62] ,\asic/lsdram/msdram/io_dmi_wr_data[61] ,\asic/lsdram/msdram/io_dmi_wr_data[60] ,\asic/lsdram/msdram/io_dmi_wr_data[59] ,\asic/lsdram/msdram/io_dmi_wr_data[58] ,\asic/lsdram/msdram/io_dmi_wr_data[57] ,\asic/lsdram/msdram/io_dmi_wr_data[56] ,\asic/lsdram/msdram/io_dmi_wr_data[55] ,\asic/lsdram/msdram/io_dmi_wr_data[54] ,\asic/lsdram/msdram/io_dmi_wr_data[53] ,\asic/lsdram/msdram/io_dmi_wr_data[52] ,\asic/lsdram/msdram/io_dmi_wr_data[51] ,\asic/lsdram/msdram/io_dmi_wr_data[50] ,\asic/lsdram/msdram/io_dmi_wr_data[49] ,\asic/lsdram/msdram/io_dmi_wr_data[48] ,\asic/lsdram/msdram/io_dmi_wr_data[47] ,\asic/lsdram/msdram/io_dmi_wr_data[46] ,\asic/lsdram/msdram/io_dmi_wr_data[45] ,\asic/lsdram/msdram/io_dmi_wr_data[44] ,\asic/lsdram/msdram/io_dmi_wr_data[43] ,\asic/lsdram/msdram/io_dmi_wr_data[42] ,\asic/lsdram/msdram/io_dmi_wr_data[41] ,\asic/lsdram/msdram/io_dmi_wr_data[40] ,\asic/lsdram/msdram/io_dmi_wr_data[39] ,\asic/lsdram/msdram/io_dmi_wr_data[38] ,\asic/lsdram/msdram/io_dmi_wr_data[37] ,\asic/lsdram/msdram/io_dmi_wr_data[36] ,\asic/lsdram/msdram/io_dmi_wr_data[35] ,\asic/lsdram/msdram/io_dmi_wr_data[34] ,\asic/lsdram/msdram/io_dmi_wr_data[33] ,\asic/lsdram/msdram/io_dmi_wr_data[32] ,\asic/lsdram/msdram/io_dmi_wr_data[31] ,\asic/lsdram/msdram/io_dmi_wr_data[30] ,\asic/lsdram/msdram/io_dmi_wr_data[29] ,\asic/lsdram/msdram/io_dmi_wr_data[28] ,\asic/lsdram/msdram/io_dmi_wr_data[27] ,\asic/lsdram/msdram/io_dmi_wr_data[26] ,\asic/lsdram/msdram/io_dmi_wr_data[25] ,\asic/lsdram/msdram/io_dmi_wr_data[24] ,\asic/lsdram/msdram/io_dmi_wr_data[23] ,\asic/lsdram/msdram/io_dmi_wr_data[22] ,\asic/lsdram/msdram/io_dmi_wr_data[21] ,\asic/lsdram/msdram/io_dmi_wr_data[20] ,\asic/lsdram/msdram/io_dmi_wr_data[19] ,\asic/lsdram/msdram/io_dmi_wr_data[18] ,\asic/lsdram/msdram/io_dmi_wr_data[17] ,\asic/lsdram/msdram/io_dmi_wr_data[16] ,\asic/lsdram/msdram/io_dmi_wr_data[15] ,\asic/lsdram/msdram/io_dmi_wr_data[14] ,\asic/lsdram/msdram/io_dmi_wr_data[13] ,\asic/lsdram/msdram/io_dmi_wr_data[12] ,\asic/lsdram/msdram/io_dmi_wr_data[11] ,\asic/lsdram/msdram/io_dmi_wr_data[10] ,\asic/lsdram/msdram/io_dmi_wr_data[9] ,\asic/lsdram/msdram/io_dmi_wr_data[8] ,\asic/lsdram/msdram/io_dmi_wr_data[7] ,\asic/lsdram/msdram/io_dmi_wr_data[6] ,\asic/lsdram/msdram/io_dmi_wr_data[5] ,\asic/lsdram/msdram/io_dmi_wr_data[4] ,\asic/lsdram/msdram/io_dmi_wr_data[3] ,\asic/lsdram/msdram/io_dmi_wr_data[2] ,\asic/lsdram/msdram/io_dmi_wr_data[1] ,\asic/lsdram/msdram/io_dmi_wr_data[0] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[31] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[30] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[29] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[28] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[27] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[26] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[25] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[24] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[23] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[22] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[21] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[20] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[19] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[18] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[17] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[16] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[15] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[14] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[13] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[12] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[11] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[10] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[9] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[8] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[7] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[6] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[5] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[4] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[3] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[2] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[1] ,\asic/lsdram/msdram/io_dmi_wr_data_mask[0] ,\asic/lsdram/msdram/io_dmi_rd_data[255] ,\asic/lsdram/msdram/io_dmi_rd_data[254] ,\asic/lsdram/msdram/io_dmi_rd_data[253] ,\asic/lsdram/msdram/io_dmi_rd_data[252] ,\asic/lsdram/msdram/io_dmi_rd_data[251] ,\asic/lsdram/msdram/io_dmi_rd_data[250] ,\asic/lsdram/msdram/io_dmi_rd_data[249] ,\asic/lsdram/msdram/io_dmi_rd_data[248] ,\asic/lsdram/msdram/io_dmi_rd_data[247] ,\asic/lsdram/msdram/io_dmi_rd_data[246] ,\asic/lsdram/msdram/io_dmi_rd_data[245] ,\asic/lsdram/msdram/io_dmi_rd_data[244] ,\asic/lsdram/msdram/io_dmi_rd_data[243] ,\asic/lsdram/msdram/io_dmi_rd_data[242] ,\asic/lsdram/msdram/io_dmi_rd_data[241] ,\asic/lsdram/msdram/io_dmi_rd_data[240] ,\asic/lsdram/msdram/io_dmi_rd_data[239] ,\asic/lsdram/msdram/io_dmi_rd_data[238] ,\asic/lsdram/msdram/io_dmi_rd_data[237] ,\asic/lsdram/msdram/io_dmi_rd_data[236] ,\asic/lsdram/msdram/io_dmi_rd_data[235] ,\asic/lsdram/msdram/io_dmi_rd_data[234] ,\asic/lsdram/msdram/io_dmi_rd_data[233] ,\asic/lsdram/msdram/io_dmi_rd_data[232] ,\asic/lsdram/msdram/io_dmi_rd_data[231] ,\asic/lsdram/msdram/io_dmi_rd_data[230] ,\asic/lsdram/msdram/io_dmi_rd_data[229] ,\asic/lsdram/msdram/io_dmi_rd_data[228] ,\asic/lsdram/msdram/io_dmi_rd_data[227] ,\asic/lsdram/msdram/io_dmi_rd_data[226] ,\asic/lsdram/msdram/io_dmi_rd_data[225] ,\asic/lsdram/msdram/io_dmi_rd_data[224] ,\asic/lsdram/msdram/io_dmi_rd_data[223] ,\asic/lsdram/msdram/io_dmi_rd_data[222] ,\asic/lsdram/msdram/io_dmi_rd_data[221] ,\asic/lsdram/msdram/io_dmi_rd_data[220] ,\asic/lsdram/msdram/io_dmi_rd_data[219] ,\asic/lsdram/msdram/io_dmi_rd_data[218] ,\asic/lsdram/msdram/io_dmi_rd_data[217] ,\asic/lsdram/msdram/io_dmi_rd_data[216] ,\asic/lsdram/msdram/io_dmi_rd_data[215] ,\asic/lsdram/msdram/io_dmi_rd_data[214] ,\asic/lsdram/msdram/io_dmi_rd_data[213] ,\asic/lsdram/msdram/io_dmi_rd_data[212] ,\asic/lsdram/msdram/io_dmi_rd_data[211] ,\asic/lsdram/msdram/io_dmi_rd_data[210] ,\asic/lsdram/msdram/io_dmi_rd_data[209] ,\asic/lsdram/msdram/io_dmi_rd_data[208] ,\asic/lsdram/msdram/io_dmi_rd_data[207] ,\asic/lsdram/msdram/io_dmi_rd_data[206] ,\asic/lsdram/msdram/io_dmi_rd_data[205] ,\asic/lsdram/msdram/io_dmi_rd_data[204] ,\asic/lsdram/msdram/io_dmi_rd_data[203] ,\asic/lsdram/msdram/io_dmi_rd_data[202] ,\asic/lsdram/msdram/io_dmi_rd_data[201] ,\asic/lsdram/msdram/io_dmi_rd_data[200] ,\asic/lsdram/msdram/io_dmi_rd_data[199] ,\asic/lsdram/msdram/io_dmi_rd_data[198] ,\asic/lsdram/msdram/io_dmi_rd_data[197] ,\asic/lsdram/msdram/io_dmi_rd_data[196] ,\asic/lsdram/msdram/io_dmi_rd_data[195] ,\asic/lsdram/msdram/io_dmi_rd_data[194] ,\asic/lsdram/msdram/io_dmi_rd_data[193] ,\asic/lsdram/msdram/io_dmi_rd_data[192] ,\asic/lsdram/msdram/io_dmi_rd_data[191] ,\asic/lsdram/msdram/io_dmi_rd_data[190] ,\asic/lsdram/msdram/io_dmi_rd_data[189] ,\asic/lsdram/msdram/io_dmi_rd_data[188] ,\asic/lsdram/msdram/io_dmi_rd_data[187] ,\asic/lsdram/msdram/io_dmi_rd_data[186] ,\asic/lsdram/msdram/io_dmi_rd_data[185] ,\asic/lsdram/msdram/io_dmi_rd_data[184] ,\asic/lsdram/msdram/io_dmi_rd_data[183] ,\asic/lsdram/msdram/io_dmi_rd_data[182] ,\asic/lsdram/msdram/io_dmi_rd_data[181] ,\asic/lsdram/msdram/io_dmi_rd_data[180] ,\asic/lsdram/msdram/io_dmi_rd_data[179] ,\asic/lsdram/msdram/io_dmi_rd_data[178] ,\asic/lsdram/msdram/io_dmi_rd_data[177] ,\asic/lsdram/msdram/io_dmi_rd_data[176] ,\asic/lsdram/msdram/io_dmi_rd_data[175] ,\asic/lsdram/msdram/io_dmi_rd_data[174] ,\asic/lsdram/msdram/io_dmi_rd_data[173] ,\asic/lsdram/msdram/io_dmi_rd_data[172] ,\asic/lsdram/msdram/io_dmi_rd_data[171] ,\asic/lsdram/msdram/io_dmi_rd_data[170] ,\asic/lsdram/msdram/io_dmi_rd_data[169] ,\asic/lsdram/msdram/io_dmi_rd_data[168] ,\asic/lsdram/msdram/io_dmi_rd_data[167] ,\asic/lsdram/msdram/io_dmi_rd_data[166] ,\asic/lsdram/msdram/io_dmi_rd_data[165] ,\asic/lsdram/msdram/io_dmi_rd_data[164] ,\asic/lsdram/msdram/io_dmi_rd_data[163] ,\asic/lsdram/msdram/io_dmi_rd_data[162] ,\asic/lsdram/msdram/io_dmi_rd_data[161] ,\asic/lsdram/msdram/io_dmi_rd_data[160] ,\asic/lsdram/msdram/io_dmi_rd_data[159] ,\asic/lsdram/msdram/io_dmi_rd_data[158] ,\asic/lsdram/msdram/io_dmi_rd_data[157] ,\asic/lsdram/msdram/io_dmi_rd_data[156] ,\asic/lsdram/msdram/io_dmi_rd_data[155] ,\asic/lsdram/msdram/io_dmi_rd_data[154] ,\asic/lsdram/msdram/io_dmi_rd_data[153] ,\asic/lsdram/msdram/io_dmi_rd_data[152] ,\asic/lsdram/msdram/io_dmi_rd_data[151] ,\asic/lsdram/msdram/io_dmi_rd_data[150] ,\asic/lsdram/msdram/io_dmi_rd_data[149] ,\asic/lsdram/msdram/io_dmi_rd_data[148] ,\asic/lsdram/msdram/io_dmi_rd_data[147] ,\asic/lsdram/msdram/io_dmi_rd_data[146] ,\asic/lsdram/msdram/io_dmi_rd_data[145] ,\asic/lsdram/msdram/io_dmi_rd_data[144] ,\asic/lsdram/msdram/io_dmi_rd_data[143] ,\asic/lsdram/msdram/io_dmi_rd_data[142] ,\asic/lsdram/msdram/io_dmi_rd_data[141] ,\asic/lsdram/msdram/io_dmi_rd_data[140] ,\asic/lsdram/msdram/io_dmi_rd_data[139] ,\asic/lsdram/msdram/io_dmi_rd_data[138] ,\asic/lsdram/msdram/io_dmi_rd_data[137] ,\asic/lsdram/msdram/io_dmi_rd_data[136] ,\asic/lsdram/msdram/io_dmi_rd_data[135] ,\asic/lsdram/msdram/io_dmi_rd_data[134] ,\asic/lsdram/msdram/io_dmi_rd_data[133] ,\asic/lsdram/msdram/io_dmi_rd_data[132] ,\asic/lsdram/msdram/io_dmi_rd_data[131] ,\asic/lsdram/msdram/io_dmi_rd_data[130] ,\asic/lsdram/msdram/io_dmi_rd_data[129] ,\asic/lsdram/msdram/io_dmi_rd_data[128] ,\asic/lsdram/msdram/io_dmi_rd_data[127] ,\asic/lsdram/msdram/io_dmi_rd_data[126] ,\asic/lsdram/msdram/io_dmi_rd_data[125] ,\asic/lsdram/msdram/io_dmi_rd_data[124] ,\asic/lsdram/msdram/io_dmi_rd_data[123] ,\asic/lsdram/msdram/io_dmi_rd_data[122] ,\asic/lsdram/msdram/io_dmi_rd_data[121] ,\asic/lsdram/msdram/io_dmi_rd_data[120] ,\asic/lsdram/msdram/io_dmi_rd_data[119] ,\asic/lsdram/msdram/io_dmi_rd_data[118] ,\asic/lsdram/msdram/io_dmi_rd_data[117] ,\asic/lsdram/msdram/io_dmi_rd_data[116] ,\asic/lsdram/msdram/io_dmi_rd_data[115] ,\asic/lsdram/msdram/io_dmi_rd_data[114] ,\asic/lsdram/msdram/io_dmi_rd_data[113] ,\asic/lsdram/msdram/io_dmi_rd_data[112] ,\asic/lsdram/msdram/io_dmi_rd_data[111] ,\asic/lsdram/msdram/io_dmi_rd_data[110] ,\asic/lsdram/msdram/io_dmi_rd_data[109] ,\asic/lsdram/msdram/io_dmi_rd_data[108] ,\asic/lsdram/msdram/io_dmi_rd_data[107] ,\asic/lsdram/msdram/io_dmi_rd_data[106] ,\asic/lsdram/msdram/io_dmi_rd_data[105] ,\asic/lsdram/msdram/io_dmi_rd_data[104] ,\asic/lsdram/msdram/io_dmi_rd_data[103] ,\asic/lsdram/msdram/io_dmi_rd_data[102] ,\asic/lsdram/msdram/io_dmi_rd_data[101] ,\asic/lsdram/msdram/io_dmi_rd_data[100] ,\asic/lsdram/msdram/io_dmi_rd_data[99] ,\asic/lsdram/msdram/io_dmi_rd_data[98] ,\asic/lsdram/msdram/io_dmi_rd_data[97] ,\asic/lsdram/msdram/io_dmi_rd_data[96] ,\asic/lsdram/msdram/io_dmi_rd_data[95] ,\asic/lsdram/msdram/io_dmi_rd_data[94] ,\asic/lsdram/msdram/io_dmi_rd_data[93] ,\asic/lsdram/msdram/io_dmi_rd_data[92] ,\asic/lsdram/msdram/io_dmi_rd_data[91] ,\asic/lsdram/msdram/io_dmi_rd_data[90] ,\asic/lsdram/msdram/io_dmi_rd_data[89] ,\asic/lsdram/msdram/io_dmi_rd_data[88] ,\asic/lsdram/msdram/io_dmi_rd_data[87] ,\asic/lsdram/msdram/io_dmi_rd_data[86] ,\asic/lsdram/msdram/io_dmi_rd_data[85] ,\asic/lsdram/msdram/io_dmi_rd_data[84] ,\asic/lsdram/msdram/io_dmi_rd_data[83] ,\asic/lsdram/msdram/io_dmi_rd_data[82] ,\asic/lsdram/msdram/io_dmi_rd_data[81] ,\asic/lsdram/msdram/io_dmi_rd_data[80] ,\asic/lsdram/msdram/io_dmi_rd_data[79] ,\asic/lsdram/msdram/io_dmi_rd_data[78] ,\asic/lsdram/msdram/io_dmi_rd_data[77] ,\asic/lsdram/msdram/io_dmi_rd_data[76] ,\asic/lsdram/msdram/io_dmi_rd_data[75] ,\asic/lsdram/msdram/io_dmi_rd_data[74] ,\asic/lsdram/msdram/io_dmi_rd_data[73] ,\asic/lsdram/msdram/io_dmi_rd_data[72] ,\asic/lsdram/msdram/io_dmi_rd_data[71] ,\asic/lsdram/msdram/io_dmi_rd_data[70] ,\asic/lsdram/msdram/io_dmi_rd_data[69] ,\asic/lsdram/msdram/io_dmi_rd_data[68] ,\asic/lsdram/msdram/io_dmi_rd_data[67] ,\asic/lsdram/msdram/io_dmi_rd_data[66] ,\asic/lsdram/msdram/io_dmi_rd_data[65] ,\asic/lsdram/msdram/io_dmi_rd_data[64] ,\asic/lsdram/msdram/io_dmi_rd_data[63] ,\asic/lsdram/msdram/io_dmi_rd_data[62] ,\asic/lsdram/msdram/io_dmi_rd_data[61] ,\asic/lsdram/msdram/io_dmi_rd_data[60] ,\asic/lsdram/msdram/io_dmi_rd_data[59] ,\asic/lsdram/msdram/io_dmi_rd_data[58] ,\asic/lsdram/msdram/io_dmi_rd_data[57] ,\asic/lsdram/msdram/io_dmi_rd_data[56] ,\asic/lsdram/msdram/io_dmi_rd_data[55] ,\asic/lsdram/msdram/io_dmi_rd_data[54] ,\asic/lsdram/msdram/io_dmi_rd_data[53] ,\asic/lsdram/msdram/io_dmi_rd_data[52] ,\asic/lsdram/msdram/io_dmi_rd_data[51] ,\asic/lsdram/msdram/io_dmi_rd_data[50] ,\asic/lsdram/msdram/io_dmi_rd_data[49] ,\asic/lsdram/msdram/io_dmi_rd_data[48] ,\asic/lsdram/msdram/io_dmi_rd_data[47] ,\asic/lsdram/msdram/io_dmi_rd_data[46] ,\asic/lsdram/msdram/io_dmi_rd_data[45] ,\asic/lsdram/msdram/io_dmi_rd_data[44] ,\asic/lsdram/msdram/io_dmi_rd_data[43] ,\asic/lsdram/msdram/io_dmi_rd_data[42] ,\asic/lsdram/msdram/io_dmi_rd_data[41] ,\asic/lsdram/msdram/io_dmi_rd_data[40] ,\asic/lsdram/msdram/io_dmi_rd_data[39] ,\asic/lsdram/msdram/io_dmi_rd_data[38] ,\asic/lsdram/msdram/io_dmi_rd_data[37] ,\asic/lsdram/msdram/io_dmi_rd_data[36] ,\asic/lsdram/msdram/io_dmi_rd_data[35] ,\asic/lsdram/msdram/io_dmi_rd_data[34] ,\asic/lsdram/msdram/io_dmi_rd_data[33] ,\asic/lsdram/msdram/io_dmi_rd_data[32] ,\asic/lsdram/msdram/io_dmi_rd_data[31] ,\asic/lsdram/msdram/io_dmi_rd_data[30] ,\asic/lsdram/msdram/io_dmi_rd_data[29] ,\asic/lsdram/msdram/io_dmi_rd_data[28] ,\asic/lsdram/msdram/io_dmi_rd_data[27] ,\asic/lsdram/msdram/io_dmi_rd_data[26] ,\asic/lsdram/msdram/io_dmi_rd_data[25] ,\asic/lsdram/msdram/io_dmi_rd_data[24] ,\asic/lsdram/msdram/io_dmi_rd_data[23] ,\asic/lsdram/msdram/io_dmi_rd_data[22] ,\asic/lsdram/msdram/io_dmi_rd_data[21] ,\asic/lsdram/msdram/io_dmi_rd_data[20] ,\asic/lsdram/msdram/io_dmi_rd_data[19] ,\asic/lsdram/msdram/io_dmi_rd_data[18] ,\asic/lsdram/msdram/io_dmi_rd_data[17] ,\asic/lsdram/msdram/io_dmi_rd_data[16] ,\asic/lsdram/msdram/io_dmi_rd_data[15] ,\asic/lsdram/msdram/io_dmi_rd_data[14] ,\asic/lsdram/msdram/io_dmi_rd_data[13] ,\asic/lsdram/msdram/io_dmi_rd_data[12] ,\asic/lsdram/msdram/io_dmi_rd_data[11] ,\asic/lsdram/msdram/io_dmi_rd_data[10] ,\asic/lsdram/msdram/io_dmi_rd_data[9] ,\asic/lsdram/msdram/io_dmi_rd_data[8] ,\asic/lsdram/msdram/io_dmi_rd_data[7] ,\asic/lsdram/msdram/io_dmi_rd_data[6] ,\asic/lsdram/msdram/io_dmi_rd_data[5] ,\asic/lsdram/msdram/io_dmi_rd_data[4] ,\asic/lsdram/msdram/io_dmi_rd_data[3] ,\asic/lsdram/msdram/io_dmi_rd_data[2] ,\asic/lsdram/msdram/io_dmi_rd_data[1] ,\asic/lsdram/msdram/io_dmi_rd_data[0] ,\asic/lsdram/msdram/io_in_rdata_r[255] ,\asic/lsdram/msdram/io_in_rdata_r[254] ,\asic/lsdram/msdram/io_in_rdata_r[253] ,\asic/lsdram/msdram/io_in_rdata_r[252] ,\asic/lsdram/msdram/io_in_rdata_r[251] ,\asic/lsdram/msdram/io_in_rdata_r[250] ,\asic/lsdram/msdram/io_in_rdata_r[249] ,\asic/lsdram/msdram/io_in_rdata_r[248] ,\asic/lsdram/msdram/io_in_rdata_r[247] ,\asic/lsdram/msdram/io_in_rdata_r[246] ,\asic/lsdram/msdram/io_in_rdata_r[245] ,\asic/lsdram/msdram/io_in_rdata_r[244] ,\asic/lsdram/msdram/io_in_rdata_r[243] ,\asic/lsdram/msdram/io_in_rdata_r[242] ,\asic/lsdram/msdram/io_in_rdata_r[241] ,\asic/lsdram/msdram/io_in_rdata_r[240] ,\asic/lsdram/msdram/io_in_rdata_r[239] ,\asic/lsdram/msdram/io_in_rdata_r[238] ,\asic/lsdram/msdram/io_in_rdata_r[237] ,\asic/lsdram/msdram/io_in_rdata_r[236] ,\asic/lsdram/msdram/io_in_rdata_r[235] ,\asic/lsdram/msdram/io_in_rdata_r[234] ,\asic/lsdram/msdram/io_in_rdata_r[233] ,\asic/lsdram/msdram/io_in_rdata_r[232] ,\asic/lsdram/msdram/io_in_rdata_r[231] ,\asic/lsdram/msdram/io_in_rdata_r[230] ,\asic/lsdram/msdram/io_in_rdata_r[229] ,\asic/lsdram/msdram/io_in_rdata_r[228] ,\asic/lsdram/msdram/io_in_rdata_r[227] ,\asic/lsdram/msdram/io_in_rdata_r[226] ,\asic/lsdram/msdram/io_in_rdata_r[225] ,\asic/lsdram/msdram/io_in_rdata_r[224] ,\asic/lsdram/msdram/io_in_rdata_r[223] ,\asic/lsdram/msdram/io_in_rdata_r[222] ,\asic/lsdram/msdram/io_in_rdata_r[221] ,\asic/lsdram/msdram/io_in_rdata_r[220] ,\asic/lsdram/msdram/io_in_rdata_r[219] ,\asic/lsdram/msdram/io_in_rdata_r[218] ,\asic/lsdram/msdram/io_in_rdata_r[217] ,\asic/lsdram/msdram/io_in_rdata_r[216] ,\asic/lsdram/msdram/io_in_rdata_r[215] ,\asic/lsdram/msdram/io_in_rdata_r[214] ,\asic/lsdram/msdram/io_in_rdata_r[213] ,\asic/lsdram/msdram/io_in_rdata_r[212] ,\asic/lsdram/msdram/io_in_rdata_r[211] ,\asic/lsdram/msdram/io_in_rdata_r[210] ,\asic/lsdram/msdram/io_in_rdata_r[209] ,\asic/lsdram/msdram/io_in_rdata_r[208] ,\asic/lsdram/msdram/io_in_rdata_r[207] ,\asic/lsdram/msdram/io_in_rdata_r[206] ,\asic/lsdram/msdram/io_in_rdata_r[205] ,\asic/lsdram/msdram/io_in_rdata_r[204] ,\asic/lsdram/msdram/io_in_rdata_r[203] ,\asic/lsdram/msdram/io_in_rdata_r[202] ,\asic/lsdram/msdram/io_in_rdata_r[201] ,\asic/lsdram/msdram/io_in_rdata_r[200] ,\asic/lsdram/msdram/io_in_rdata_r[199] ,\asic/lsdram/msdram/io_in_rdata_r[198] ,\asic/lsdram/msdram/io_in_rdata_r[197] ,\asic/lsdram/msdram/io_in_rdata_r[196] ,\asic/lsdram/msdram/io_in_rdata_r[195] ,\asic/lsdram/msdram/io_in_rdata_r[194] ,\asic/lsdram/msdram/io_in_rdata_r[193] ,\asic/lsdram/msdram/io_in_rdata_r[192] ,\asic/lsdram/msdram/io_in_rdata_r[191] ,\asic/lsdram/msdram/io_in_rdata_r[190] ,\asic/lsdram/msdram/io_in_rdata_r[189] ,\asic/lsdram/msdram/io_in_rdata_r[188] ,\asic/lsdram/msdram/io_in_rdata_r[187] ,\asic/lsdram/msdram/io_in_rdata_r[186] ,\asic/lsdram/msdram/io_in_rdata_r[185] ,\asic/lsdram/msdram/io_in_rdata_r[184] ,\asic/lsdram/msdram/io_in_rdata_r[183] ,\asic/lsdram/msdram/io_in_rdata_r[182] ,\asic/lsdram/msdram/io_in_rdata_r[181] ,\asic/lsdram/msdram/io_in_rdata_r[180] ,\asic/lsdram/msdram/io_in_rdata_r[179] ,\asic/lsdram/msdram/io_in_rdata_r[178] ,\asic/lsdram/msdram/io_in_rdata_r[177] ,\asic/lsdram/msdram/io_in_rdata_r[176] ,\asic/lsdram/msdram/io_in_rdata_r[175] ,\asic/lsdram/msdram/io_in_rdata_r[174] ,\asic/lsdram/msdram/io_in_rdata_r[173] ,\asic/lsdram/msdram/io_in_rdata_r[172] ,\asic/lsdram/msdram/io_in_rdata_r[171] ,\asic/lsdram/msdram/io_in_rdata_r[170] ,\asic/lsdram/msdram/io_in_rdata_r[169] ,\asic/lsdram/msdram/io_in_rdata_r[168] ,\asic/lsdram/msdram/io_in_rdata_r[167] ,\asic/lsdram/msdram/io_in_rdata_r[166] ,\asic/lsdram/msdram/io_in_rdata_r[165] ,\asic/lsdram/msdram/io_in_rdata_r[164] ,\asic/lsdram/msdram/io_in_rdata_r[163] ,\asic/lsdram/msdram/io_in_rdata_r[162] ,\asic/lsdram/msdram/io_in_rdata_r[161] ,\asic/lsdram/msdram/io_in_rdata_r[160] ,\asic/lsdram/msdram/io_in_rdata_r[159] ,\asic/lsdram/msdram/io_in_rdata_r[158] ,\asic/lsdram/msdram/io_in_rdata_r[157] ,\asic/lsdram/msdram/io_in_rdata_r[156] ,\asic/lsdram/msdram/io_in_rdata_r[155] ,\asic/lsdram/msdram/io_in_rdata_r[154] ,\asic/lsdram/msdram/io_in_rdata_r[153] ,\asic/lsdram/msdram/io_in_rdata_r[152] ,\asic/lsdram/msdram/io_in_rdata_r[151] ,\asic/lsdram/msdram/io_in_rdata_r[150] ,\asic/lsdram/msdram/io_in_rdata_r[149] ,\asic/lsdram/msdram/io_in_rdata_r[148] ,\asic/lsdram/msdram/io_in_rdata_r[147] ,\asic/lsdram/msdram/io_in_rdata_r[146] ,\asic/lsdram/msdram/io_in_rdata_r[145] ,\asic/lsdram/msdram/io_in_rdata_r[144] ,\asic/lsdram/msdram/io_in_rdata_r[143] ,\asic/lsdram/msdram/io_in_rdata_r[142] ,\asic/lsdram/msdram/io_in_rdata_r[141] ,\asic/lsdram/msdram/io_in_rdata_r[140] ,\asic/lsdram/msdram/io_in_rdata_r[139] ,\asic/lsdram/msdram/io_in_rdata_r[138] ,\asic/lsdram/msdram/io_in_rdata_r[137] ,\asic/lsdram/msdram/io_in_rdata_r[136] ,\asic/lsdram/msdram/io_in_rdata_r[135] ,\asic/lsdram/msdram/io_in_rdata_r[134] ,\asic/lsdram/msdram/io_in_rdata_r[133] ,\asic/lsdram/msdram/io_in_rdata_r[132] ,\asic/lsdram/msdram/io_in_rdata_r[131] ,\asic/lsdram/msdram/io_in_rdata_r[130] ,\asic/lsdram/msdram/io_in_rdata_r[129] ,\asic/lsdram/msdram/io_in_rdata_r[128] ,\asic/lsdram/msdram/io_in_rdata_r[127] ,\asic/lsdram/msdram/io_in_rdata_r[126] ,\asic/lsdram/msdram/io_in_rdata_r[125] ,\asic/lsdram/msdram/io_in_rdata_r[124] ,\asic/lsdram/msdram/io_in_rdata_r[123] ,\asic/lsdram/msdram/io_in_rdata_r[122] ,\asic/lsdram/msdram/io_in_rdata_r[121] ,\asic/lsdram/msdram/io_in_rdata_r[120] ,\asic/lsdram/msdram/io_in_rdata_r[119] ,\asic/lsdram/msdram/io_in_rdata_r[118] ,\asic/lsdram/msdram/io_in_rdata_r[117] ,\asic/lsdram/msdram/io_in_rdata_r[116] ,\asic/lsdram/msdram/io_in_rdata_r[115] ,\asic/lsdram/msdram/io_in_rdata_r[114] ,\asic/lsdram/msdram/io_in_rdata_r[113] ,\asic/lsdram/msdram/io_in_rdata_r[112] ,\asic/lsdram/msdram/io_in_rdata_r[111] ,\asic/lsdram/msdram/io_in_rdata_r[110] ,\asic/lsdram/msdram/io_in_rdata_r[109] ,\asic/lsdram/msdram/io_in_rdata_r[108] ,\asic/lsdram/msdram/io_in_rdata_r[107] ,\asic/lsdram/msdram/io_in_rdata_r[106] ,\asic/lsdram/msdram/io_in_rdata_r[105] ,\asic/lsdram/msdram/io_in_rdata_r[104] ,\asic/lsdram/msdram/io_in_rdata_r[103] ,\asic/lsdram/msdram/io_in_rdata_r[102] ,\asic/lsdram/msdram/io_in_rdata_r[101] ,\asic/lsdram/msdram/io_in_rdata_r[100] ,\asic/lsdram/msdram/io_in_rdata_r[99] ,\asic/lsdram/msdram/io_in_rdata_r[98] ,\asic/lsdram/msdram/io_in_rdata_r[97] ,\asic/lsdram/msdram/io_in_rdata_r[96] ,\asic/lsdram/msdram/io_in_rdata_r[95] ,\asic/lsdram/msdram/io_in_rdata_r[94] ,\asic/lsdram/msdram/io_in_rdata_r[93] ,\asic/lsdram/msdram/io_in_rdata_r[92] ,\asic/lsdram/msdram/io_in_rdata_r[91] ,\asic/lsdram/msdram/io_in_rdata_r[90] ,\asic/lsdram/msdram/io_in_rdata_r[89] ,\asic/lsdram/msdram/io_in_rdata_r[88] ,\asic/lsdram/msdram/io_in_rdata_r[87] ,\asic/lsdram/msdram/io_in_rdata_r[86] ,\asic/lsdram/msdram/io_in_rdata_r[85] ,\asic/lsdram/msdram/io_in_rdata_r[84] ,\asic/lsdram/msdram/io_in_rdata_r[83] ,\asic/lsdram/msdram/io_in_rdata_r[82] ,\asic/lsdram/msdram/io_in_rdata_r[81] ,\asic/lsdram/msdram/io_in_rdata_r[80] ,\asic/lsdram/msdram/io_in_rdata_r[79] ,\asic/lsdram/msdram/io_in_rdata_r[78] ,\asic/lsdram/msdram/io_in_rdata_r[77] ,\asic/lsdram/msdram/io_in_rdata_r[76] ,\asic/lsdram/msdram/io_in_rdata_r[75] ,\asic/lsdram/msdram/io_in_rdata_r[74] ,\asic/lsdram/msdram/io_in_rdata_r[73] ,\asic/lsdram/msdram/io_in_rdata_r[72] ,\asic/lsdram/msdram/io_in_rdata_r[71] ,\asic/lsdram/msdram/io_in_rdata_r[70] ,\asic/lsdram/msdram/io_in_rdata_r[69] ,\asic/lsdram/msdram/io_in_rdata_r[68] ,\asic/lsdram/msdram/io_in_rdata_r[67] ,\asic/lsdram/msdram/io_in_rdata_r[66] ,\asic/lsdram/msdram/io_in_rdata_r[65] ,\asic/lsdram/msdram/io_in_rdata_r[64] ,\asic/lsdram/msdram/io_in_rdata_r[63] ,\asic/lsdram/msdram/io_in_rdata_r[62] ,\asic/lsdram/msdram/io_in_rdata_r[61] ,\asic/lsdram/msdram/io_in_rdata_r[60] ,\asic/lsdram/msdram/io_in_rdata_r[59] ,\asic/lsdram/msdram/io_in_rdata_r[58] ,\asic/lsdram/msdram/io_in_rdata_r[57] ,\asic/lsdram/msdram/io_in_rdata_r[56] ,\asic/lsdram/msdram/io_in_rdata_r[55] ,\asic/lsdram/msdram/io_in_rdata_r[54] ,\asic/lsdram/msdram/io_in_rdata_r[53] ,\asic/lsdram/msdram/io_in_rdata_r[52] ,\asic/lsdram/msdram/io_in_rdata_r[51] ,\asic/lsdram/msdram/io_in_rdata_r[50] ,\asic/lsdram/msdram/io_in_rdata_r[49] ,\asic/lsdram/msdram/io_in_rdata_r[48] ,\asic/lsdram/msdram/io_in_rdata_r[47] ,\asic/lsdram/msdram/io_in_rdata_r[46] ,\asic/lsdram/msdram/io_in_rdata_r[45] ,\asic/lsdram/msdram/io_in_rdata_r[44] ,\asic/lsdram/msdram/io_in_rdata_r[43] ,\asic/lsdram/msdram/io_in_rdata_r[42] ,\asic/lsdram/msdram/io_in_rdata_r[41] ,\asic/lsdram/msdram/io_in_rdata_r[40] ,\asic/lsdram/msdram/io_in_rdata_r[39] ,\asic/lsdram/msdram/io_in_rdata_r[38] ,\asic/lsdram/msdram/io_in_rdata_r[37] ,\asic/lsdram/msdram/io_in_rdata_r[36] ,\asic/lsdram/msdram/io_in_rdata_r[35] ,\asic/lsdram/msdram/io_in_rdata_r[34] ,\asic/lsdram/msdram/io_in_rdata_r[33] ,\asic/lsdram/msdram/io_in_rdata_r[32] ,\asic/lsdram/msdram/io_in_rdata_r[31] ,\asic/lsdram/msdram/io_in_rdata_r[30] ,\asic/lsdram/msdram/io_in_rdata_r[29] ,\asic/lsdram/msdram/io_in_rdata_r[28] ,\asic/lsdram/msdram/io_in_rdata_r[27] ,\asic/lsdram/msdram/io_in_rdata_r[26] ,\asic/lsdram/msdram/io_in_rdata_r[25] ,\asic/lsdram/msdram/io_in_rdata_r[24] ,\asic/lsdram/msdram/io_in_rdata_r[23] ,\asic/lsdram/msdram/io_in_rdata_r[22] ,\asic/lsdram/msdram/io_in_rdata_r[21] ,\asic/lsdram/msdram/io_in_rdata_r[20] ,\asic/lsdram/msdram/io_in_rdata_r[19] ,\asic/lsdram/msdram/io_in_rdata_r[18] ,\asic/lsdram/msdram/io_in_rdata_r[17] ,\asic/lsdram/msdram/io_in_rdata_r[16] ,\asic/lsdram/msdram/io_in_rdata_r[15] ,\asic/lsdram/msdram/io_in_rdata_r[14] ,\asic/lsdram/msdram/io_in_rdata_r[13] ,\asic/lsdram/msdram/io_in_rdata_r[12] ,\asic/lsdram/msdram/io_in_rdata_r[11] ,\asic/lsdram/msdram/io_in_rdata_r[10] ,\asic/lsdram/msdram/io_in_rdata_r[9] ,\asic/lsdram/msdram/io_in_rdata_r[8] ,\asic/lsdram/msdram/io_in_rdata_r[7] ,\asic/lsdram/msdram/io_in_rdata_r[6] ,\asic/lsdram/msdram/io_in_rdata_r[5] ,\asic/lsdram/msdram/io_in_rdata_r[4] ,\asic/lsdram/msdram/io_in_rdata_r[3] ,\asic/lsdram/msdram/io_in_rdata_r[2] ,\asic/lsdram/msdram/io_in_rdata_r[1] ,\asic/lsdram/msdram/io_in_rdata_r[0] ,\asic/lsdram/msdram/io_clk_out ,\asic/lsdram/msdram/io_in_awready ,\asic/lsdram/msdram/io_in_awvalid ,\asic/lsdram/msdram/io_in_wready ,\asic/lsdram/msdram/io_in_wvalid ,\asic/lsdram/msdram/io_in_bready ,\asic/lsdram/msdram/io_in_bvalid ,\asic/lsdram/msdram/io_in_arready ,\asic/lsdram/msdram/io_in_arvalid ,\asic/lsdram/msdram/io_in_rready ,\asic/lsdram/msdram/io_in_rvalid ,\asic/lsdram/msdram/io_dmi_cmd_en ,\asic/lsdram/msdram/io_dmi_wr_data_en ,\asic/lsdram/msdram/io_dmi_wr_data_end ,\asic/lsdram/msdram/io_dmi_clk_out ,\asic/lsdram/msdram/io_dmi_init_calib_complete ,\asic/lsdram/msdram/io_dmi_cmd_ready ,\asic/lsdram/msdram/io_dmi_wr_data_rdy ,\asic/lsdram/msdram/io_dmi_rd_data_valid }),
    .clk_i(clock)
);

endmodule
