//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03
//Part Number: GW5AST-LV138FPG676AC2/I1
//Device: GW5AST-138B
//Device Version: B
//Created Time: Sat May 18 21:02:03 2024

module SRAM_SDPB (dout, clka, cea, clkb, ceb, oce, reset, ada, din, adb, byte_ena);

output [31:0] dout;
input clka;
input cea;
input clkb;
input ceb;
input oce;
input reset;
input [16:0] ada;
input [31:0] din;
input [16:0] adb;
input [3:0] byte_ena;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire lut_f_64;
wire lut_f_65;
wire lut_f_66;
wire lut_f_67;
wire lut_f_68;
wire lut_f_69;
wire lut_f_70;
wire lut_f_71;
wire lut_f_72;
wire lut_f_73;
wire lut_f_74;
wire lut_f_75;
wire lut_f_76;
wire lut_f_77;
wire lut_f_78;
wire lut_f_79;
wire lut_f_80;
wire lut_f_81;
wire lut_f_82;
wire lut_f_83;
wire lut_f_84;
wire lut_f_85;
wire lut_f_86;
wire lut_f_87;
wire lut_f_88;
wire lut_f_89;
wire lut_f_90;
wire lut_f_91;
wire lut_f_92;
wire lut_f_93;
wire lut_f_94;
wire lut_f_95;
wire lut_f_96;
wire lut_f_97;
wire lut_f_98;
wire lut_f_99;
wire lut_f_100;
wire lut_f_101;
wire lut_f_102;
wire lut_f_103;
wire lut_f_104;
wire lut_f_105;
wire lut_f_106;
wire lut_f_107;
wire lut_f_108;
wire lut_f_109;
wire lut_f_110;
wire lut_f_111;
wire lut_f_112;
wire lut_f_113;
wire lut_f_114;
wire lut_f_115;
wire lut_f_116;
wire lut_f_117;
wire lut_f_118;
wire lut_f_119;
wire lut_f_120;
wire lut_f_121;
wire lut_f_122;
wire lut_f_123;
wire lut_f_124;
wire lut_f_125;
wire lut_f_126;
wire lut_f_127;
wire lut_f_128;
wire lut_f_129;
wire lut_f_130;
wire lut_f_131;
wire lut_f_132;
wire lut_f_133;
wire lut_f_134;
wire lut_f_135;
wire lut_f_136;
wire lut_f_137;
wire lut_f_138;
wire lut_f_139;
wire lut_f_140;
wire lut_f_141;
wire lut_f_142;
wire lut_f_143;
wire lut_f_144;
wire lut_f_145;
wire lut_f_146;
wire lut_f_147;
wire lut_f_148;
wire lut_f_149;
wire lut_f_150;
wire lut_f_151;
wire lut_f_152;
wire lut_f_153;
wire lut_f_154;
wire lut_f_155;
wire lut_f_156;
wire lut_f_157;
wire lut_f_158;
wire lut_f_159;
wire lut_f_160;
wire lut_f_161;
wire lut_f_162;
wire lut_f_163;
wire lut_f_164;
wire lut_f_165;
wire lut_f_166;
wire lut_f_167;
wire lut_f_168;
wire lut_f_169;
wire lut_f_170;
wire lut_f_171;
wire lut_f_172;
wire lut_f_173;
wire lut_f_174;
wire lut_f_175;
wire lut_f_176;
wire lut_f_177;
wire lut_f_178;
wire lut_f_179;
wire lut_f_180;
wire lut_f_181;
wire lut_f_182;
wire lut_f_183;
wire lut_f_184;
wire lut_f_185;
wire lut_f_186;
wire lut_f_187;
wire lut_f_188;
wire lut_f_189;
wire lut_f_190;
wire lut_f_191;
wire lut_f_192;
wire lut_f_193;
wire lut_f_194;
wire lut_f_195;
wire lut_f_196;
wire lut_f_197;
wire lut_f_198;
wire lut_f_199;
wire lut_f_200;
wire lut_f_201;
wire lut_f_202;
wire lut_f_203;
wire lut_f_204;
wire lut_f_205;
wire lut_f_206;
wire lut_f_207;
wire lut_f_208;
wire lut_f_209;
wire lut_f_210;
wire lut_f_211;
wire lut_f_212;
wire lut_f_213;
wire lut_f_214;
wire lut_f_215;
wire lut_f_216;
wire lut_f_217;
wire lut_f_218;
wire lut_f_219;
wire lut_f_220;
wire lut_f_221;
wire lut_f_222;
wire lut_f_223;
wire lut_f_224;
wire lut_f_225;
wire lut_f_226;
wire lut_f_227;
wire lut_f_228;
wire lut_f_229;
wire lut_f_230;
wire lut_f_231;
wire lut_f_232;
wire lut_f_233;
wire lut_f_234;
wire lut_f_235;
wire lut_f_236;
wire lut_f_237;
wire lut_f_238;
wire lut_f_239;
wire lut_f_240;
wire lut_f_241;
wire lut_f_242;
wire lut_f_243;
wire lut_f_244;
wire lut_f_245;
wire lut_f_246;
wire lut_f_247;
wire lut_f_248;
wire lut_f_249;
wire lut_f_250;
wire lut_f_251;
wire lut_f_252;
wire lut_f_253;
wire lut_f_254;
wire lut_f_255;
wire [15:0] sdpb_inst_0_dout_w;
wire [15:0] sdpb_inst_0_dout;
wire [15:0] sdpb_inst_1_dout_w;
wire [15:0] sdpb_inst_1_dout;
wire [15:0] sdpb_inst_2_dout_w;
wire [15:0] sdpb_inst_2_dout;
wire [15:0] sdpb_inst_3_dout_w;
wire [15:0] sdpb_inst_3_dout;
wire [15:0] sdpb_inst_4_dout_w;
wire [15:0] sdpb_inst_4_dout;
wire [15:0] sdpb_inst_5_dout_w;
wire [15:0] sdpb_inst_5_dout;
wire [15:0] sdpb_inst_6_dout_w;
wire [15:0] sdpb_inst_6_dout;
wire [15:0] sdpb_inst_7_dout_w;
wire [15:0] sdpb_inst_7_dout;
wire [15:0] sdpb_inst_8_dout_w;
wire [15:0] sdpb_inst_8_dout;
wire [15:0] sdpb_inst_9_dout_w;
wire [15:0] sdpb_inst_9_dout;
wire [15:0] sdpb_inst_10_dout_w;
wire [15:0] sdpb_inst_10_dout;
wire [15:0] sdpb_inst_11_dout_w;
wire [15:0] sdpb_inst_11_dout;
wire [15:0] sdpb_inst_12_dout_w;
wire [15:0] sdpb_inst_12_dout;
wire [15:0] sdpb_inst_13_dout_w;
wire [15:0] sdpb_inst_13_dout;
wire [15:0] sdpb_inst_14_dout_w;
wire [15:0] sdpb_inst_14_dout;
wire [15:0] sdpb_inst_15_dout_w;
wire [15:0] sdpb_inst_15_dout;
wire [15:0] sdpb_inst_16_dout_w;
wire [15:0] sdpb_inst_16_dout;
wire [15:0] sdpb_inst_17_dout_w;
wire [15:0] sdpb_inst_17_dout;
wire [15:0] sdpb_inst_18_dout_w;
wire [15:0] sdpb_inst_18_dout;
wire [15:0] sdpb_inst_19_dout_w;
wire [15:0] sdpb_inst_19_dout;
wire [15:0] sdpb_inst_20_dout_w;
wire [15:0] sdpb_inst_20_dout;
wire [15:0] sdpb_inst_21_dout_w;
wire [15:0] sdpb_inst_21_dout;
wire [15:0] sdpb_inst_22_dout_w;
wire [15:0] sdpb_inst_22_dout;
wire [15:0] sdpb_inst_23_dout_w;
wire [15:0] sdpb_inst_23_dout;
wire [15:0] sdpb_inst_24_dout_w;
wire [15:0] sdpb_inst_24_dout;
wire [15:0] sdpb_inst_25_dout_w;
wire [15:0] sdpb_inst_25_dout;
wire [15:0] sdpb_inst_26_dout_w;
wire [15:0] sdpb_inst_26_dout;
wire [15:0] sdpb_inst_27_dout_w;
wire [15:0] sdpb_inst_27_dout;
wire [15:0] sdpb_inst_28_dout_w;
wire [15:0] sdpb_inst_28_dout;
wire [15:0] sdpb_inst_29_dout_w;
wire [15:0] sdpb_inst_29_dout;
wire [15:0] sdpb_inst_30_dout_w;
wire [15:0] sdpb_inst_30_dout;
wire [15:0] sdpb_inst_31_dout_w;
wire [15:0] sdpb_inst_31_dout;
wire [15:0] sdpb_inst_32_dout_w;
wire [15:0] sdpb_inst_32_dout;
wire [15:0] sdpb_inst_33_dout_w;
wire [15:0] sdpb_inst_33_dout;
wire [15:0] sdpb_inst_34_dout_w;
wire [15:0] sdpb_inst_34_dout;
wire [15:0] sdpb_inst_35_dout_w;
wire [15:0] sdpb_inst_35_dout;
wire [15:0] sdpb_inst_36_dout_w;
wire [15:0] sdpb_inst_36_dout;
wire [15:0] sdpb_inst_37_dout_w;
wire [15:0] sdpb_inst_37_dout;
wire [15:0] sdpb_inst_38_dout_w;
wire [15:0] sdpb_inst_38_dout;
wire [15:0] sdpb_inst_39_dout_w;
wire [15:0] sdpb_inst_39_dout;
wire [15:0] sdpb_inst_40_dout_w;
wire [15:0] sdpb_inst_40_dout;
wire [15:0] sdpb_inst_41_dout_w;
wire [15:0] sdpb_inst_41_dout;
wire [15:0] sdpb_inst_42_dout_w;
wire [15:0] sdpb_inst_42_dout;
wire [15:0] sdpb_inst_43_dout_w;
wire [15:0] sdpb_inst_43_dout;
wire [15:0] sdpb_inst_44_dout_w;
wire [15:0] sdpb_inst_44_dout;
wire [15:0] sdpb_inst_45_dout_w;
wire [15:0] sdpb_inst_45_dout;
wire [15:0] sdpb_inst_46_dout_w;
wire [15:0] sdpb_inst_46_dout;
wire [15:0] sdpb_inst_47_dout_w;
wire [15:0] sdpb_inst_47_dout;
wire [15:0] sdpb_inst_48_dout_w;
wire [15:0] sdpb_inst_48_dout;
wire [15:0] sdpb_inst_49_dout_w;
wire [15:0] sdpb_inst_49_dout;
wire [15:0] sdpb_inst_50_dout_w;
wire [15:0] sdpb_inst_50_dout;
wire [15:0] sdpb_inst_51_dout_w;
wire [15:0] sdpb_inst_51_dout;
wire [15:0] sdpb_inst_52_dout_w;
wire [15:0] sdpb_inst_52_dout;
wire [15:0] sdpb_inst_53_dout_w;
wire [15:0] sdpb_inst_53_dout;
wire [15:0] sdpb_inst_54_dout_w;
wire [15:0] sdpb_inst_54_dout;
wire [15:0] sdpb_inst_55_dout_w;
wire [15:0] sdpb_inst_55_dout;
wire [15:0] sdpb_inst_56_dout_w;
wire [15:0] sdpb_inst_56_dout;
wire [15:0] sdpb_inst_57_dout_w;
wire [15:0] sdpb_inst_57_dout;
wire [15:0] sdpb_inst_58_dout_w;
wire [15:0] sdpb_inst_58_dout;
wire [15:0] sdpb_inst_59_dout_w;
wire [15:0] sdpb_inst_59_dout;
wire [15:0] sdpb_inst_60_dout_w;
wire [15:0] sdpb_inst_60_dout;
wire [15:0] sdpb_inst_61_dout_w;
wire [15:0] sdpb_inst_61_dout;
wire [15:0] sdpb_inst_62_dout_w;
wire [15:0] sdpb_inst_62_dout;
wire [15:0] sdpb_inst_63_dout_w;
wire [15:0] sdpb_inst_63_dout;
wire [15:0] sdpb_inst_64_dout_w;
wire [15:0] sdpb_inst_64_dout;
wire [15:0] sdpb_inst_65_dout_w;
wire [15:0] sdpb_inst_65_dout;
wire [15:0] sdpb_inst_66_dout_w;
wire [15:0] sdpb_inst_66_dout;
wire [15:0] sdpb_inst_67_dout_w;
wire [15:0] sdpb_inst_67_dout;
wire [15:0] sdpb_inst_68_dout_w;
wire [15:0] sdpb_inst_68_dout;
wire [15:0] sdpb_inst_69_dout_w;
wire [15:0] sdpb_inst_69_dout;
wire [15:0] sdpb_inst_70_dout_w;
wire [15:0] sdpb_inst_70_dout;
wire [15:0] sdpb_inst_71_dout_w;
wire [15:0] sdpb_inst_71_dout;
wire [15:0] sdpb_inst_72_dout_w;
wire [15:0] sdpb_inst_72_dout;
wire [15:0] sdpb_inst_73_dout_w;
wire [15:0] sdpb_inst_73_dout;
wire [15:0] sdpb_inst_74_dout_w;
wire [15:0] sdpb_inst_74_dout;
wire [15:0] sdpb_inst_75_dout_w;
wire [15:0] sdpb_inst_75_dout;
wire [15:0] sdpb_inst_76_dout_w;
wire [15:0] sdpb_inst_76_dout;
wire [15:0] sdpb_inst_77_dout_w;
wire [15:0] sdpb_inst_77_dout;
wire [15:0] sdpb_inst_78_dout_w;
wire [15:0] sdpb_inst_78_dout;
wire [15:0] sdpb_inst_79_dout_w;
wire [15:0] sdpb_inst_79_dout;
wire [15:0] sdpb_inst_80_dout_w;
wire [15:0] sdpb_inst_80_dout;
wire [15:0] sdpb_inst_81_dout_w;
wire [15:0] sdpb_inst_81_dout;
wire [15:0] sdpb_inst_82_dout_w;
wire [15:0] sdpb_inst_82_dout;
wire [15:0] sdpb_inst_83_dout_w;
wire [15:0] sdpb_inst_83_dout;
wire [15:0] sdpb_inst_84_dout_w;
wire [15:0] sdpb_inst_84_dout;
wire [15:0] sdpb_inst_85_dout_w;
wire [15:0] sdpb_inst_85_dout;
wire [15:0] sdpb_inst_86_dout_w;
wire [15:0] sdpb_inst_86_dout;
wire [15:0] sdpb_inst_87_dout_w;
wire [15:0] sdpb_inst_87_dout;
wire [15:0] sdpb_inst_88_dout_w;
wire [15:0] sdpb_inst_88_dout;
wire [15:0] sdpb_inst_89_dout_w;
wire [15:0] sdpb_inst_89_dout;
wire [15:0] sdpb_inst_90_dout_w;
wire [15:0] sdpb_inst_90_dout;
wire [15:0] sdpb_inst_91_dout_w;
wire [15:0] sdpb_inst_91_dout;
wire [15:0] sdpb_inst_92_dout_w;
wire [15:0] sdpb_inst_92_dout;
wire [15:0] sdpb_inst_93_dout_w;
wire [15:0] sdpb_inst_93_dout;
wire [15:0] sdpb_inst_94_dout_w;
wire [15:0] sdpb_inst_94_dout;
wire [15:0] sdpb_inst_95_dout_w;
wire [15:0] sdpb_inst_95_dout;
wire [15:0] sdpb_inst_96_dout_w;
wire [15:0] sdpb_inst_96_dout;
wire [15:0] sdpb_inst_97_dout_w;
wire [15:0] sdpb_inst_97_dout;
wire [15:0] sdpb_inst_98_dout_w;
wire [15:0] sdpb_inst_98_dout;
wire [15:0] sdpb_inst_99_dout_w;
wire [15:0] sdpb_inst_99_dout;
wire [15:0] sdpb_inst_100_dout_w;
wire [15:0] sdpb_inst_100_dout;
wire [15:0] sdpb_inst_101_dout_w;
wire [15:0] sdpb_inst_101_dout;
wire [15:0] sdpb_inst_102_dout_w;
wire [15:0] sdpb_inst_102_dout;
wire [15:0] sdpb_inst_103_dout_w;
wire [15:0] sdpb_inst_103_dout;
wire [15:0] sdpb_inst_104_dout_w;
wire [15:0] sdpb_inst_104_dout;
wire [15:0] sdpb_inst_105_dout_w;
wire [15:0] sdpb_inst_105_dout;
wire [15:0] sdpb_inst_106_dout_w;
wire [15:0] sdpb_inst_106_dout;
wire [15:0] sdpb_inst_107_dout_w;
wire [15:0] sdpb_inst_107_dout;
wire [15:0] sdpb_inst_108_dout_w;
wire [15:0] sdpb_inst_108_dout;
wire [15:0] sdpb_inst_109_dout_w;
wire [15:0] sdpb_inst_109_dout;
wire [15:0] sdpb_inst_110_dout_w;
wire [15:0] sdpb_inst_110_dout;
wire [15:0] sdpb_inst_111_dout_w;
wire [15:0] sdpb_inst_111_dout;
wire [15:0] sdpb_inst_112_dout_w;
wire [15:0] sdpb_inst_112_dout;
wire [15:0] sdpb_inst_113_dout_w;
wire [15:0] sdpb_inst_113_dout;
wire [15:0] sdpb_inst_114_dout_w;
wire [15:0] sdpb_inst_114_dout;
wire [15:0] sdpb_inst_115_dout_w;
wire [15:0] sdpb_inst_115_dout;
wire [15:0] sdpb_inst_116_dout_w;
wire [15:0] sdpb_inst_116_dout;
wire [15:0] sdpb_inst_117_dout_w;
wire [15:0] sdpb_inst_117_dout;
wire [15:0] sdpb_inst_118_dout_w;
wire [15:0] sdpb_inst_118_dout;
wire [15:0] sdpb_inst_119_dout_w;
wire [15:0] sdpb_inst_119_dout;
wire [15:0] sdpb_inst_120_dout_w;
wire [15:0] sdpb_inst_120_dout;
wire [15:0] sdpb_inst_121_dout_w;
wire [15:0] sdpb_inst_121_dout;
wire [15:0] sdpb_inst_122_dout_w;
wire [15:0] sdpb_inst_122_dout;
wire [15:0] sdpb_inst_123_dout_w;
wire [15:0] sdpb_inst_123_dout;
wire [15:0] sdpb_inst_124_dout_w;
wire [15:0] sdpb_inst_124_dout;
wire [15:0] sdpb_inst_125_dout_w;
wire [15:0] sdpb_inst_125_dout;
wire [15:0] sdpb_inst_126_dout_w;
wire [15:0] sdpb_inst_126_dout;
wire [15:0] sdpb_inst_127_dout_w;
wire [15:0] sdpb_inst_127_dout;
wire [15:0] sdpb_inst_128_dout_w;
wire [31:16] sdpb_inst_128_dout;
wire [15:0] sdpb_inst_129_dout_w;
wire [31:16] sdpb_inst_129_dout;
wire [15:0] sdpb_inst_130_dout_w;
wire [31:16] sdpb_inst_130_dout;
wire [15:0] sdpb_inst_131_dout_w;
wire [31:16] sdpb_inst_131_dout;
wire [15:0] sdpb_inst_132_dout_w;
wire [31:16] sdpb_inst_132_dout;
wire [15:0] sdpb_inst_133_dout_w;
wire [31:16] sdpb_inst_133_dout;
wire [15:0] sdpb_inst_134_dout_w;
wire [31:16] sdpb_inst_134_dout;
wire [15:0] sdpb_inst_135_dout_w;
wire [31:16] sdpb_inst_135_dout;
wire [15:0] sdpb_inst_136_dout_w;
wire [31:16] sdpb_inst_136_dout;
wire [15:0] sdpb_inst_137_dout_w;
wire [31:16] sdpb_inst_137_dout;
wire [15:0] sdpb_inst_138_dout_w;
wire [31:16] sdpb_inst_138_dout;
wire [15:0] sdpb_inst_139_dout_w;
wire [31:16] sdpb_inst_139_dout;
wire [15:0] sdpb_inst_140_dout_w;
wire [31:16] sdpb_inst_140_dout;
wire [15:0] sdpb_inst_141_dout_w;
wire [31:16] sdpb_inst_141_dout;
wire [15:0] sdpb_inst_142_dout_w;
wire [31:16] sdpb_inst_142_dout;
wire [15:0] sdpb_inst_143_dout_w;
wire [31:16] sdpb_inst_143_dout;
wire [15:0] sdpb_inst_144_dout_w;
wire [31:16] sdpb_inst_144_dout;
wire [15:0] sdpb_inst_145_dout_w;
wire [31:16] sdpb_inst_145_dout;
wire [15:0] sdpb_inst_146_dout_w;
wire [31:16] sdpb_inst_146_dout;
wire [15:0] sdpb_inst_147_dout_w;
wire [31:16] sdpb_inst_147_dout;
wire [15:0] sdpb_inst_148_dout_w;
wire [31:16] sdpb_inst_148_dout;
wire [15:0] sdpb_inst_149_dout_w;
wire [31:16] sdpb_inst_149_dout;
wire [15:0] sdpb_inst_150_dout_w;
wire [31:16] sdpb_inst_150_dout;
wire [15:0] sdpb_inst_151_dout_w;
wire [31:16] sdpb_inst_151_dout;
wire [15:0] sdpb_inst_152_dout_w;
wire [31:16] sdpb_inst_152_dout;
wire [15:0] sdpb_inst_153_dout_w;
wire [31:16] sdpb_inst_153_dout;
wire [15:0] sdpb_inst_154_dout_w;
wire [31:16] sdpb_inst_154_dout;
wire [15:0] sdpb_inst_155_dout_w;
wire [31:16] sdpb_inst_155_dout;
wire [15:0] sdpb_inst_156_dout_w;
wire [31:16] sdpb_inst_156_dout;
wire [15:0] sdpb_inst_157_dout_w;
wire [31:16] sdpb_inst_157_dout;
wire [15:0] sdpb_inst_158_dout_w;
wire [31:16] sdpb_inst_158_dout;
wire [15:0] sdpb_inst_159_dout_w;
wire [31:16] sdpb_inst_159_dout;
wire [15:0] sdpb_inst_160_dout_w;
wire [31:16] sdpb_inst_160_dout;
wire [15:0] sdpb_inst_161_dout_w;
wire [31:16] sdpb_inst_161_dout;
wire [15:0] sdpb_inst_162_dout_w;
wire [31:16] sdpb_inst_162_dout;
wire [15:0] sdpb_inst_163_dout_w;
wire [31:16] sdpb_inst_163_dout;
wire [15:0] sdpb_inst_164_dout_w;
wire [31:16] sdpb_inst_164_dout;
wire [15:0] sdpb_inst_165_dout_w;
wire [31:16] sdpb_inst_165_dout;
wire [15:0] sdpb_inst_166_dout_w;
wire [31:16] sdpb_inst_166_dout;
wire [15:0] sdpb_inst_167_dout_w;
wire [31:16] sdpb_inst_167_dout;
wire [15:0] sdpb_inst_168_dout_w;
wire [31:16] sdpb_inst_168_dout;
wire [15:0] sdpb_inst_169_dout_w;
wire [31:16] sdpb_inst_169_dout;
wire [15:0] sdpb_inst_170_dout_w;
wire [31:16] sdpb_inst_170_dout;
wire [15:0] sdpb_inst_171_dout_w;
wire [31:16] sdpb_inst_171_dout;
wire [15:0] sdpb_inst_172_dout_w;
wire [31:16] sdpb_inst_172_dout;
wire [15:0] sdpb_inst_173_dout_w;
wire [31:16] sdpb_inst_173_dout;
wire [15:0] sdpb_inst_174_dout_w;
wire [31:16] sdpb_inst_174_dout;
wire [15:0] sdpb_inst_175_dout_w;
wire [31:16] sdpb_inst_175_dout;
wire [15:0] sdpb_inst_176_dout_w;
wire [31:16] sdpb_inst_176_dout;
wire [15:0] sdpb_inst_177_dout_w;
wire [31:16] sdpb_inst_177_dout;
wire [15:0] sdpb_inst_178_dout_w;
wire [31:16] sdpb_inst_178_dout;
wire [15:0] sdpb_inst_179_dout_w;
wire [31:16] sdpb_inst_179_dout;
wire [15:0] sdpb_inst_180_dout_w;
wire [31:16] sdpb_inst_180_dout;
wire [15:0] sdpb_inst_181_dout_w;
wire [31:16] sdpb_inst_181_dout;
wire [15:0] sdpb_inst_182_dout_w;
wire [31:16] sdpb_inst_182_dout;
wire [15:0] sdpb_inst_183_dout_w;
wire [31:16] sdpb_inst_183_dout;
wire [15:0] sdpb_inst_184_dout_w;
wire [31:16] sdpb_inst_184_dout;
wire [15:0] sdpb_inst_185_dout_w;
wire [31:16] sdpb_inst_185_dout;
wire [15:0] sdpb_inst_186_dout_w;
wire [31:16] sdpb_inst_186_dout;
wire [15:0] sdpb_inst_187_dout_w;
wire [31:16] sdpb_inst_187_dout;
wire [15:0] sdpb_inst_188_dout_w;
wire [31:16] sdpb_inst_188_dout;
wire [15:0] sdpb_inst_189_dout_w;
wire [31:16] sdpb_inst_189_dout;
wire [15:0] sdpb_inst_190_dout_w;
wire [31:16] sdpb_inst_190_dout;
wire [15:0] sdpb_inst_191_dout_w;
wire [31:16] sdpb_inst_191_dout;
wire [15:0] sdpb_inst_192_dout_w;
wire [31:16] sdpb_inst_192_dout;
wire [15:0] sdpb_inst_193_dout_w;
wire [31:16] sdpb_inst_193_dout;
wire [15:0] sdpb_inst_194_dout_w;
wire [31:16] sdpb_inst_194_dout;
wire [15:0] sdpb_inst_195_dout_w;
wire [31:16] sdpb_inst_195_dout;
wire [15:0] sdpb_inst_196_dout_w;
wire [31:16] sdpb_inst_196_dout;
wire [15:0] sdpb_inst_197_dout_w;
wire [31:16] sdpb_inst_197_dout;
wire [15:0] sdpb_inst_198_dout_w;
wire [31:16] sdpb_inst_198_dout;
wire [15:0] sdpb_inst_199_dout_w;
wire [31:16] sdpb_inst_199_dout;
wire [15:0] sdpb_inst_200_dout_w;
wire [31:16] sdpb_inst_200_dout;
wire [15:0] sdpb_inst_201_dout_w;
wire [31:16] sdpb_inst_201_dout;
wire [15:0] sdpb_inst_202_dout_w;
wire [31:16] sdpb_inst_202_dout;
wire [15:0] sdpb_inst_203_dout_w;
wire [31:16] sdpb_inst_203_dout;
wire [15:0] sdpb_inst_204_dout_w;
wire [31:16] sdpb_inst_204_dout;
wire [15:0] sdpb_inst_205_dout_w;
wire [31:16] sdpb_inst_205_dout;
wire [15:0] sdpb_inst_206_dout_w;
wire [31:16] sdpb_inst_206_dout;
wire [15:0] sdpb_inst_207_dout_w;
wire [31:16] sdpb_inst_207_dout;
wire [15:0] sdpb_inst_208_dout_w;
wire [31:16] sdpb_inst_208_dout;
wire [15:0] sdpb_inst_209_dout_w;
wire [31:16] sdpb_inst_209_dout;
wire [15:0] sdpb_inst_210_dout_w;
wire [31:16] sdpb_inst_210_dout;
wire [15:0] sdpb_inst_211_dout_w;
wire [31:16] sdpb_inst_211_dout;
wire [15:0] sdpb_inst_212_dout_w;
wire [31:16] sdpb_inst_212_dout;
wire [15:0] sdpb_inst_213_dout_w;
wire [31:16] sdpb_inst_213_dout;
wire [15:0] sdpb_inst_214_dout_w;
wire [31:16] sdpb_inst_214_dout;
wire [15:0] sdpb_inst_215_dout_w;
wire [31:16] sdpb_inst_215_dout;
wire [15:0] sdpb_inst_216_dout_w;
wire [31:16] sdpb_inst_216_dout;
wire [15:0] sdpb_inst_217_dout_w;
wire [31:16] sdpb_inst_217_dout;
wire [15:0] sdpb_inst_218_dout_w;
wire [31:16] sdpb_inst_218_dout;
wire [15:0] sdpb_inst_219_dout_w;
wire [31:16] sdpb_inst_219_dout;
wire [15:0] sdpb_inst_220_dout_w;
wire [31:16] sdpb_inst_220_dout;
wire [15:0] sdpb_inst_221_dout_w;
wire [31:16] sdpb_inst_221_dout;
wire [15:0] sdpb_inst_222_dout_w;
wire [31:16] sdpb_inst_222_dout;
wire [15:0] sdpb_inst_223_dout_w;
wire [31:16] sdpb_inst_223_dout;
wire [15:0] sdpb_inst_224_dout_w;
wire [31:16] sdpb_inst_224_dout;
wire [15:0] sdpb_inst_225_dout_w;
wire [31:16] sdpb_inst_225_dout;
wire [15:0] sdpb_inst_226_dout_w;
wire [31:16] sdpb_inst_226_dout;
wire [15:0] sdpb_inst_227_dout_w;
wire [31:16] sdpb_inst_227_dout;
wire [15:0] sdpb_inst_228_dout_w;
wire [31:16] sdpb_inst_228_dout;
wire [15:0] sdpb_inst_229_dout_w;
wire [31:16] sdpb_inst_229_dout;
wire [15:0] sdpb_inst_230_dout_w;
wire [31:16] sdpb_inst_230_dout;
wire [15:0] sdpb_inst_231_dout_w;
wire [31:16] sdpb_inst_231_dout;
wire [15:0] sdpb_inst_232_dout_w;
wire [31:16] sdpb_inst_232_dout;
wire [15:0] sdpb_inst_233_dout_w;
wire [31:16] sdpb_inst_233_dout;
wire [15:0] sdpb_inst_234_dout_w;
wire [31:16] sdpb_inst_234_dout;
wire [15:0] sdpb_inst_235_dout_w;
wire [31:16] sdpb_inst_235_dout;
wire [15:0] sdpb_inst_236_dout_w;
wire [31:16] sdpb_inst_236_dout;
wire [15:0] sdpb_inst_237_dout_w;
wire [31:16] sdpb_inst_237_dout;
wire [15:0] sdpb_inst_238_dout_w;
wire [31:16] sdpb_inst_238_dout;
wire [15:0] sdpb_inst_239_dout_w;
wire [31:16] sdpb_inst_239_dout;
wire [15:0] sdpb_inst_240_dout_w;
wire [31:16] sdpb_inst_240_dout;
wire [15:0] sdpb_inst_241_dout_w;
wire [31:16] sdpb_inst_241_dout;
wire [15:0] sdpb_inst_242_dout_w;
wire [31:16] sdpb_inst_242_dout;
wire [15:0] sdpb_inst_243_dout_w;
wire [31:16] sdpb_inst_243_dout;
wire [15:0] sdpb_inst_244_dout_w;
wire [31:16] sdpb_inst_244_dout;
wire [15:0] sdpb_inst_245_dout_w;
wire [31:16] sdpb_inst_245_dout;
wire [15:0] sdpb_inst_246_dout_w;
wire [31:16] sdpb_inst_246_dout;
wire [15:0] sdpb_inst_247_dout_w;
wire [31:16] sdpb_inst_247_dout;
wire [15:0] sdpb_inst_248_dout_w;
wire [31:16] sdpb_inst_248_dout;
wire [15:0] sdpb_inst_249_dout_w;
wire [31:16] sdpb_inst_249_dout;
wire [15:0] sdpb_inst_250_dout_w;
wire [31:16] sdpb_inst_250_dout;
wire [15:0] sdpb_inst_251_dout_w;
wire [31:16] sdpb_inst_251_dout;
wire [15:0] sdpb_inst_252_dout_w;
wire [31:16] sdpb_inst_252_dout;
wire [15:0] sdpb_inst_253_dout_w;
wire [31:16] sdpb_inst_253_dout;
wire [15:0] sdpb_inst_254_dout_w;
wire [31:16] sdpb_inst_254_dout;
wire [15:0] sdpb_inst_255_dout_w;
wire [31:16] sdpb_inst_255_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_503;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_588;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_629;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_755;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_867;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_881;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_898;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_929;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_944;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_960;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire mux_o_991;
wire mux_o_992;
wire mux_o_993;
wire mux_o_994;
wire mux_o_995;
wire mux_o_996;
wire mux_o_997;
wire mux_o_998;
wire mux_o_999;
wire mux_o_1000;
wire mux_o_1001;
wire mux_o_1002;
wire mux_o_1003;
wire mux_o_1004;
wire mux_o_1005;
wire mux_o_1006;
wire mux_o_1007;
wire mux_o_1008;
wire mux_o_1009;
wire mux_o_1010;
wire mux_o_1011;
wire mux_o_1012;
wire mux_o_1013;
wire mux_o_1014;
wire mux_o_1016;
wire mux_o_1017;
wire mux_o_1018;
wire mux_o_1019;
wire mux_o_1020;
wire mux_o_1021;
wire mux_o_1022;
wire mux_o_1023;
wire mux_o_1024;
wire mux_o_1025;
wire mux_o_1026;
wire mux_o_1027;
wire mux_o_1028;
wire mux_o_1029;
wire mux_o_1030;
wire mux_o_1031;
wire mux_o_1032;
wire mux_o_1033;
wire mux_o_1034;
wire mux_o_1035;
wire mux_o_1036;
wire mux_o_1037;
wire mux_o_1038;
wire mux_o_1039;
wire mux_o_1040;
wire mux_o_1041;
wire mux_o_1042;
wire mux_o_1043;
wire mux_o_1044;
wire mux_o_1045;
wire mux_o_1046;
wire mux_o_1047;
wire mux_o_1048;
wire mux_o_1049;
wire mux_o_1050;
wire mux_o_1051;
wire mux_o_1052;
wire mux_o_1053;
wire mux_o_1054;
wire mux_o_1055;
wire mux_o_1056;
wire mux_o_1057;
wire mux_o_1058;
wire mux_o_1059;
wire mux_o_1060;
wire mux_o_1061;
wire mux_o_1062;
wire mux_o_1063;
wire mux_o_1064;
wire mux_o_1065;
wire mux_o_1066;
wire mux_o_1067;
wire mux_o_1068;
wire mux_o_1069;
wire mux_o_1070;
wire mux_o_1071;
wire mux_o_1072;
wire mux_o_1073;
wire mux_o_1074;
wire mux_o_1075;
wire mux_o_1076;
wire mux_o_1077;
wire mux_o_1078;
wire mux_o_1079;
wire mux_o_1080;
wire mux_o_1081;
wire mux_o_1082;
wire mux_o_1083;
wire mux_o_1084;
wire mux_o_1085;
wire mux_o_1086;
wire mux_o_1087;
wire mux_o_1088;
wire mux_o_1089;
wire mux_o_1090;
wire mux_o_1091;
wire mux_o_1092;
wire mux_o_1093;
wire mux_o_1094;
wire mux_o_1095;
wire mux_o_1096;
wire mux_o_1097;
wire mux_o_1098;
wire mux_o_1099;
wire mux_o_1100;
wire mux_o_1101;
wire mux_o_1102;
wire mux_o_1103;
wire mux_o_1104;
wire mux_o_1105;
wire mux_o_1106;
wire mux_o_1107;
wire mux_o_1108;
wire mux_o_1109;
wire mux_o_1110;
wire mux_o_1111;
wire mux_o_1112;
wire mux_o_1113;
wire mux_o_1114;
wire mux_o_1115;
wire mux_o_1116;
wire mux_o_1117;
wire mux_o_1118;
wire mux_o_1119;
wire mux_o_1120;
wire mux_o_1121;
wire mux_o_1122;
wire mux_o_1123;
wire mux_o_1124;
wire mux_o_1125;
wire mux_o_1126;
wire mux_o_1127;
wire mux_o_1128;
wire mux_o_1129;
wire mux_o_1130;
wire mux_o_1131;
wire mux_o_1132;
wire mux_o_1133;
wire mux_o_1134;
wire mux_o_1135;
wire mux_o_1136;
wire mux_o_1137;
wire mux_o_1138;
wire mux_o_1139;
wire mux_o_1140;
wire mux_o_1141;
wire mux_o_1143;
wire mux_o_1144;
wire mux_o_1145;
wire mux_o_1146;
wire mux_o_1147;
wire mux_o_1148;
wire mux_o_1149;
wire mux_o_1150;
wire mux_o_1151;
wire mux_o_1152;
wire mux_o_1153;
wire mux_o_1154;
wire mux_o_1155;
wire mux_o_1156;
wire mux_o_1157;
wire mux_o_1158;
wire mux_o_1159;
wire mux_o_1160;
wire mux_o_1161;
wire mux_o_1162;
wire mux_o_1163;
wire mux_o_1164;
wire mux_o_1165;
wire mux_o_1166;
wire mux_o_1167;
wire mux_o_1168;
wire mux_o_1169;
wire mux_o_1170;
wire mux_o_1171;
wire mux_o_1172;
wire mux_o_1173;
wire mux_o_1174;
wire mux_o_1175;
wire mux_o_1176;
wire mux_o_1177;
wire mux_o_1178;
wire mux_o_1179;
wire mux_o_1180;
wire mux_o_1181;
wire mux_o_1182;
wire mux_o_1183;
wire mux_o_1184;
wire mux_o_1185;
wire mux_o_1186;
wire mux_o_1187;
wire mux_o_1188;
wire mux_o_1189;
wire mux_o_1190;
wire mux_o_1191;
wire mux_o_1192;
wire mux_o_1193;
wire mux_o_1194;
wire mux_o_1195;
wire mux_o_1196;
wire mux_o_1197;
wire mux_o_1198;
wire mux_o_1199;
wire mux_o_1200;
wire mux_o_1201;
wire mux_o_1202;
wire mux_o_1203;
wire mux_o_1204;
wire mux_o_1205;
wire mux_o_1206;
wire mux_o_1207;
wire mux_o_1208;
wire mux_o_1209;
wire mux_o_1210;
wire mux_o_1211;
wire mux_o_1212;
wire mux_o_1213;
wire mux_o_1214;
wire mux_o_1215;
wire mux_o_1216;
wire mux_o_1217;
wire mux_o_1218;
wire mux_o_1219;
wire mux_o_1220;
wire mux_o_1221;
wire mux_o_1222;
wire mux_o_1223;
wire mux_o_1224;
wire mux_o_1225;
wire mux_o_1226;
wire mux_o_1227;
wire mux_o_1228;
wire mux_o_1229;
wire mux_o_1230;
wire mux_o_1231;
wire mux_o_1232;
wire mux_o_1233;
wire mux_o_1234;
wire mux_o_1235;
wire mux_o_1236;
wire mux_o_1237;
wire mux_o_1238;
wire mux_o_1239;
wire mux_o_1240;
wire mux_o_1241;
wire mux_o_1242;
wire mux_o_1243;
wire mux_o_1244;
wire mux_o_1245;
wire mux_o_1246;
wire mux_o_1247;
wire mux_o_1248;
wire mux_o_1249;
wire mux_o_1250;
wire mux_o_1251;
wire mux_o_1252;
wire mux_o_1253;
wire mux_o_1254;
wire mux_o_1255;
wire mux_o_1256;
wire mux_o_1257;
wire mux_o_1258;
wire mux_o_1259;
wire mux_o_1260;
wire mux_o_1261;
wire mux_o_1262;
wire mux_o_1263;
wire mux_o_1264;
wire mux_o_1265;
wire mux_o_1266;
wire mux_o_1267;
wire mux_o_1268;
wire mux_o_1270;
wire mux_o_1271;
wire mux_o_1272;
wire mux_o_1273;
wire mux_o_1274;
wire mux_o_1275;
wire mux_o_1276;
wire mux_o_1277;
wire mux_o_1278;
wire mux_o_1279;
wire mux_o_1280;
wire mux_o_1281;
wire mux_o_1282;
wire mux_o_1283;
wire mux_o_1284;
wire mux_o_1285;
wire mux_o_1286;
wire mux_o_1287;
wire mux_o_1288;
wire mux_o_1289;
wire mux_o_1290;
wire mux_o_1291;
wire mux_o_1292;
wire mux_o_1293;
wire mux_o_1294;
wire mux_o_1295;
wire mux_o_1296;
wire mux_o_1297;
wire mux_o_1298;
wire mux_o_1299;
wire mux_o_1300;
wire mux_o_1301;
wire mux_o_1302;
wire mux_o_1303;
wire mux_o_1304;
wire mux_o_1305;
wire mux_o_1306;
wire mux_o_1307;
wire mux_o_1308;
wire mux_o_1309;
wire mux_o_1310;
wire mux_o_1311;
wire mux_o_1312;
wire mux_o_1313;
wire mux_o_1314;
wire mux_o_1315;
wire mux_o_1316;
wire mux_o_1317;
wire mux_o_1318;
wire mux_o_1319;
wire mux_o_1320;
wire mux_o_1321;
wire mux_o_1322;
wire mux_o_1323;
wire mux_o_1324;
wire mux_o_1325;
wire mux_o_1326;
wire mux_o_1327;
wire mux_o_1328;
wire mux_o_1329;
wire mux_o_1330;
wire mux_o_1331;
wire mux_o_1332;
wire mux_o_1333;
wire mux_o_1334;
wire mux_o_1335;
wire mux_o_1336;
wire mux_o_1337;
wire mux_o_1338;
wire mux_o_1339;
wire mux_o_1340;
wire mux_o_1341;
wire mux_o_1342;
wire mux_o_1343;
wire mux_o_1344;
wire mux_o_1345;
wire mux_o_1346;
wire mux_o_1347;
wire mux_o_1348;
wire mux_o_1349;
wire mux_o_1350;
wire mux_o_1351;
wire mux_o_1352;
wire mux_o_1353;
wire mux_o_1354;
wire mux_o_1355;
wire mux_o_1356;
wire mux_o_1357;
wire mux_o_1358;
wire mux_o_1359;
wire mux_o_1360;
wire mux_o_1361;
wire mux_o_1362;
wire mux_o_1363;
wire mux_o_1364;
wire mux_o_1365;
wire mux_o_1366;
wire mux_o_1367;
wire mux_o_1368;
wire mux_o_1369;
wire mux_o_1370;
wire mux_o_1371;
wire mux_o_1372;
wire mux_o_1373;
wire mux_o_1374;
wire mux_o_1375;
wire mux_o_1376;
wire mux_o_1377;
wire mux_o_1378;
wire mux_o_1379;
wire mux_o_1380;
wire mux_o_1381;
wire mux_o_1382;
wire mux_o_1383;
wire mux_o_1384;
wire mux_o_1385;
wire mux_o_1386;
wire mux_o_1387;
wire mux_o_1388;
wire mux_o_1389;
wire mux_o_1390;
wire mux_o_1391;
wire mux_o_1392;
wire mux_o_1393;
wire mux_o_1394;
wire mux_o_1395;
wire mux_o_1397;
wire mux_o_1398;
wire mux_o_1399;
wire mux_o_1400;
wire mux_o_1401;
wire mux_o_1402;
wire mux_o_1403;
wire mux_o_1404;
wire mux_o_1405;
wire mux_o_1406;
wire mux_o_1407;
wire mux_o_1408;
wire mux_o_1409;
wire mux_o_1410;
wire mux_o_1411;
wire mux_o_1412;
wire mux_o_1413;
wire mux_o_1414;
wire mux_o_1415;
wire mux_o_1416;
wire mux_o_1417;
wire mux_o_1418;
wire mux_o_1419;
wire mux_o_1420;
wire mux_o_1421;
wire mux_o_1422;
wire mux_o_1423;
wire mux_o_1424;
wire mux_o_1425;
wire mux_o_1426;
wire mux_o_1427;
wire mux_o_1428;
wire mux_o_1429;
wire mux_o_1430;
wire mux_o_1431;
wire mux_o_1432;
wire mux_o_1433;
wire mux_o_1434;
wire mux_o_1435;
wire mux_o_1436;
wire mux_o_1437;
wire mux_o_1438;
wire mux_o_1439;
wire mux_o_1440;
wire mux_o_1441;
wire mux_o_1442;
wire mux_o_1443;
wire mux_o_1444;
wire mux_o_1445;
wire mux_o_1446;
wire mux_o_1447;
wire mux_o_1448;
wire mux_o_1449;
wire mux_o_1450;
wire mux_o_1451;
wire mux_o_1452;
wire mux_o_1453;
wire mux_o_1454;
wire mux_o_1455;
wire mux_o_1456;
wire mux_o_1457;
wire mux_o_1458;
wire mux_o_1459;
wire mux_o_1460;
wire mux_o_1461;
wire mux_o_1462;
wire mux_o_1463;
wire mux_o_1464;
wire mux_o_1465;
wire mux_o_1466;
wire mux_o_1467;
wire mux_o_1468;
wire mux_o_1469;
wire mux_o_1470;
wire mux_o_1471;
wire mux_o_1472;
wire mux_o_1473;
wire mux_o_1474;
wire mux_o_1475;
wire mux_o_1476;
wire mux_o_1477;
wire mux_o_1478;
wire mux_o_1479;
wire mux_o_1480;
wire mux_o_1481;
wire mux_o_1482;
wire mux_o_1483;
wire mux_o_1484;
wire mux_o_1485;
wire mux_o_1486;
wire mux_o_1487;
wire mux_o_1488;
wire mux_o_1489;
wire mux_o_1490;
wire mux_o_1491;
wire mux_o_1492;
wire mux_o_1493;
wire mux_o_1494;
wire mux_o_1495;
wire mux_o_1496;
wire mux_o_1497;
wire mux_o_1498;
wire mux_o_1499;
wire mux_o_1500;
wire mux_o_1501;
wire mux_o_1502;
wire mux_o_1503;
wire mux_o_1504;
wire mux_o_1505;
wire mux_o_1506;
wire mux_o_1507;
wire mux_o_1508;
wire mux_o_1509;
wire mux_o_1510;
wire mux_o_1511;
wire mux_o_1512;
wire mux_o_1513;
wire mux_o_1514;
wire mux_o_1515;
wire mux_o_1516;
wire mux_o_1517;
wire mux_o_1518;
wire mux_o_1519;
wire mux_o_1520;
wire mux_o_1521;
wire mux_o_1522;
wire mux_o_1524;
wire mux_o_1525;
wire mux_o_1526;
wire mux_o_1527;
wire mux_o_1528;
wire mux_o_1529;
wire mux_o_1530;
wire mux_o_1531;
wire mux_o_1532;
wire mux_o_1533;
wire mux_o_1534;
wire mux_o_1535;
wire mux_o_1536;
wire mux_o_1537;
wire mux_o_1538;
wire mux_o_1539;
wire mux_o_1540;
wire mux_o_1541;
wire mux_o_1542;
wire mux_o_1543;
wire mux_o_1544;
wire mux_o_1545;
wire mux_o_1546;
wire mux_o_1547;
wire mux_o_1548;
wire mux_o_1549;
wire mux_o_1550;
wire mux_o_1551;
wire mux_o_1552;
wire mux_o_1553;
wire mux_o_1554;
wire mux_o_1555;
wire mux_o_1556;
wire mux_o_1557;
wire mux_o_1558;
wire mux_o_1559;
wire mux_o_1560;
wire mux_o_1561;
wire mux_o_1562;
wire mux_o_1563;
wire mux_o_1564;
wire mux_o_1565;
wire mux_o_1566;
wire mux_o_1567;
wire mux_o_1568;
wire mux_o_1569;
wire mux_o_1570;
wire mux_o_1571;
wire mux_o_1572;
wire mux_o_1573;
wire mux_o_1574;
wire mux_o_1575;
wire mux_o_1576;
wire mux_o_1577;
wire mux_o_1578;
wire mux_o_1579;
wire mux_o_1580;
wire mux_o_1581;
wire mux_o_1582;
wire mux_o_1583;
wire mux_o_1584;
wire mux_o_1585;
wire mux_o_1586;
wire mux_o_1587;
wire mux_o_1588;
wire mux_o_1589;
wire mux_o_1590;
wire mux_o_1591;
wire mux_o_1592;
wire mux_o_1593;
wire mux_o_1594;
wire mux_o_1595;
wire mux_o_1596;
wire mux_o_1597;
wire mux_o_1598;
wire mux_o_1599;
wire mux_o_1600;
wire mux_o_1601;
wire mux_o_1602;
wire mux_o_1603;
wire mux_o_1604;
wire mux_o_1605;
wire mux_o_1606;
wire mux_o_1607;
wire mux_o_1608;
wire mux_o_1609;
wire mux_o_1610;
wire mux_o_1611;
wire mux_o_1612;
wire mux_o_1613;
wire mux_o_1614;
wire mux_o_1615;
wire mux_o_1616;
wire mux_o_1617;
wire mux_o_1618;
wire mux_o_1619;
wire mux_o_1620;
wire mux_o_1621;
wire mux_o_1622;
wire mux_o_1623;
wire mux_o_1624;
wire mux_o_1625;
wire mux_o_1626;
wire mux_o_1627;
wire mux_o_1628;
wire mux_o_1629;
wire mux_o_1630;
wire mux_o_1631;
wire mux_o_1632;
wire mux_o_1633;
wire mux_o_1634;
wire mux_o_1635;
wire mux_o_1636;
wire mux_o_1637;
wire mux_o_1638;
wire mux_o_1639;
wire mux_o_1640;
wire mux_o_1641;
wire mux_o_1642;
wire mux_o_1643;
wire mux_o_1644;
wire mux_o_1645;
wire mux_o_1646;
wire mux_o_1647;
wire mux_o_1648;
wire mux_o_1649;
wire mux_o_1651;
wire mux_o_1652;
wire mux_o_1653;
wire mux_o_1654;
wire mux_o_1655;
wire mux_o_1656;
wire mux_o_1657;
wire mux_o_1658;
wire mux_o_1659;
wire mux_o_1660;
wire mux_o_1661;
wire mux_o_1662;
wire mux_o_1663;
wire mux_o_1664;
wire mux_o_1665;
wire mux_o_1666;
wire mux_o_1667;
wire mux_o_1668;
wire mux_o_1669;
wire mux_o_1670;
wire mux_o_1671;
wire mux_o_1672;
wire mux_o_1673;
wire mux_o_1674;
wire mux_o_1675;
wire mux_o_1676;
wire mux_o_1677;
wire mux_o_1678;
wire mux_o_1679;
wire mux_o_1680;
wire mux_o_1681;
wire mux_o_1682;
wire mux_o_1683;
wire mux_o_1684;
wire mux_o_1685;
wire mux_o_1686;
wire mux_o_1687;
wire mux_o_1688;
wire mux_o_1689;
wire mux_o_1690;
wire mux_o_1691;
wire mux_o_1692;
wire mux_o_1693;
wire mux_o_1694;
wire mux_o_1695;
wire mux_o_1696;
wire mux_o_1697;
wire mux_o_1698;
wire mux_o_1699;
wire mux_o_1700;
wire mux_o_1701;
wire mux_o_1702;
wire mux_o_1703;
wire mux_o_1704;
wire mux_o_1705;
wire mux_o_1706;
wire mux_o_1707;
wire mux_o_1708;
wire mux_o_1709;
wire mux_o_1710;
wire mux_o_1711;
wire mux_o_1712;
wire mux_o_1713;
wire mux_o_1714;
wire mux_o_1715;
wire mux_o_1716;
wire mux_o_1717;
wire mux_o_1718;
wire mux_o_1719;
wire mux_o_1720;
wire mux_o_1721;
wire mux_o_1722;
wire mux_o_1723;
wire mux_o_1724;
wire mux_o_1725;
wire mux_o_1726;
wire mux_o_1727;
wire mux_o_1728;
wire mux_o_1729;
wire mux_o_1730;
wire mux_o_1731;
wire mux_o_1732;
wire mux_o_1733;
wire mux_o_1734;
wire mux_o_1735;
wire mux_o_1736;
wire mux_o_1737;
wire mux_o_1738;
wire mux_o_1739;
wire mux_o_1740;
wire mux_o_1741;
wire mux_o_1742;
wire mux_o_1743;
wire mux_o_1744;
wire mux_o_1745;
wire mux_o_1746;
wire mux_o_1747;
wire mux_o_1748;
wire mux_o_1749;
wire mux_o_1750;
wire mux_o_1751;
wire mux_o_1752;
wire mux_o_1753;
wire mux_o_1754;
wire mux_o_1755;
wire mux_o_1756;
wire mux_o_1757;
wire mux_o_1758;
wire mux_o_1759;
wire mux_o_1760;
wire mux_o_1761;
wire mux_o_1762;
wire mux_o_1763;
wire mux_o_1764;
wire mux_o_1765;
wire mux_o_1766;
wire mux_o_1767;
wire mux_o_1768;
wire mux_o_1769;
wire mux_o_1770;
wire mux_o_1771;
wire mux_o_1772;
wire mux_o_1773;
wire mux_o_1774;
wire mux_o_1775;
wire mux_o_1776;
wire mux_o_1778;
wire mux_o_1779;
wire mux_o_1780;
wire mux_o_1781;
wire mux_o_1782;
wire mux_o_1783;
wire mux_o_1784;
wire mux_o_1785;
wire mux_o_1786;
wire mux_o_1787;
wire mux_o_1788;
wire mux_o_1789;
wire mux_o_1790;
wire mux_o_1791;
wire mux_o_1792;
wire mux_o_1793;
wire mux_o_1794;
wire mux_o_1795;
wire mux_o_1796;
wire mux_o_1797;
wire mux_o_1798;
wire mux_o_1799;
wire mux_o_1800;
wire mux_o_1801;
wire mux_o_1802;
wire mux_o_1803;
wire mux_o_1804;
wire mux_o_1805;
wire mux_o_1806;
wire mux_o_1807;
wire mux_o_1808;
wire mux_o_1809;
wire mux_o_1810;
wire mux_o_1811;
wire mux_o_1812;
wire mux_o_1813;
wire mux_o_1814;
wire mux_o_1815;
wire mux_o_1816;
wire mux_o_1817;
wire mux_o_1818;
wire mux_o_1819;
wire mux_o_1820;
wire mux_o_1821;
wire mux_o_1822;
wire mux_o_1823;
wire mux_o_1824;
wire mux_o_1825;
wire mux_o_1826;
wire mux_o_1827;
wire mux_o_1828;
wire mux_o_1829;
wire mux_o_1830;
wire mux_o_1831;
wire mux_o_1832;
wire mux_o_1833;
wire mux_o_1834;
wire mux_o_1835;
wire mux_o_1836;
wire mux_o_1837;
wire mux_o_1838;
wire mux_o_1839;
wire mux_o_1840;
wire mux_o_1841;
wire mux_o_1842;
wire mux_o_1843;
wire mux_o_1844;
wire mux_o_1845;
wire mux_o_1846;
wire mux_o_1847;
wire mux_o_1848;
wire mux_o_1849;
wire mux_o_1850;
wire mux_o_1851;
wire mux_o_1852;
wire mux_o_1853;
wire mux_o_1854;
wire mux_o_1855;
wire mux_o_1856;
wire mux_o_1857;
wire mux_o_1858;
wire mux_o_1859;
wire mux_o_1860;
wire mux_o_1861;
wire mux_o_1862;
wire mux_o_1863;
wire mux_o_1864;
wire mux_o_1865;
wire mux_o_1866;
wire mux_o_1867;
wire mux_o_1868;
wire mux_o_1869;
wire mux_o_1870;
wire mux_o_1871;
wire mux_o_1872;
wire mux_o_1873;
wire mux_o_1874;
wire mux_o_1875;
wire mux_o_1876;
wire mux_o_1877;
wire mux_o_1878;
wire mux_o_1879;
wire mux_o_1880;
wire mux_o_1881;
wire mux_o_1882;
wire mux_o_1883;
wire mux_o_1884;
wire mux_o_1885;
wire mux_o_1886;
wire mux_o_1887;
wire mux_o_1888;
wire mux_o_1889;
wire mux_o_1890;
wire mux_o_1891;
wire mux_o_1892;
wire mux_o_1893;
wire mux_o_1894;
wire mux_o_1895;
wire mux_o_1896;
wire mux_o_1897;
wire mux_o_1898;
wire mux_o_1899;
wire mux_o_1900;
wire mux_o_1901;
wire mux_o_1902;
wire mux_o_1903;
wire mux_o_1905;
wire mux_o_1906;
wire mux_o_1907;
wire mux_o_1908;
wire mux_o_1909;
wire mux_o_1910;
wire mux_o_1911;
wire mux_o_1912;
wire mux_o_1913;
wire mux_o_1914;
wire mux_o_1915;
wire mux_o_1916;
wire mux_o_1917;
wire mux_o_1918;
wire mux_o_1919;
wire mux_o_1920;
wire mux_o_1921;
wire mux_o_1922;
wire mux_o_1923;
wire mux_o_1924;
wire mux_o_1925;
wire mux_o_1926;
wire mux_o_1927;
wire mux_o_1928;
wire mux_o_1929;
wire mux_o_1930;
wire mux_o_1931;
wire mux_o_1932;
wire mux_o_1933;
wire mux_o_1934;
wire mux_o_1935;
wire mux_o_1936;
wire mux_o_1937;
wire mux_o_1938;
wire mux_o_1939;
wire mux_o_1940;
wire mux_o_1941;
wire mux_o_1942;
wire mux_o_1943;
wire mux_o_1944;
wire mux_o_1945;
wire mux_o_1946;
wire mux_o_1947;
wire mux_o_1948;
wire mux_o_1949;
wire mux_o_1950;
wire mux_o_1951;
wire mux_o_1952;
wire mux_o_1953;
wire mux_o_1954;
wire mux_o_1955;
wire mux_o_1956;
wire mux_o_1957;
wire mux_o_1958;
wire mux_o_1959;
wire mux_o_1960;
wire mux_o_1961;
wire mux_o_1962;
wire mux_o_1963;
wire mux_o_1964;
wire mux_o_1965;
wire mux_o_1966;
wire mux_o_1967;
wire mux_o_1968;
wire mux_o_1969;
wire mux_o_1970;
wire mux_o_1971;
wire mux_o_1972;
wire mux_o_1973;
wire mux_o_1974;
wire mux_o_1975;
wire mux_o_1976;
wire mux_o_1977;
wire mux_o_1978;
wire mux_o_1979;
wire mux_o_1980;
wire mux_o_1981;
wire mux_o_1982;
wire mux_o_1983;
wire mux_o_1984;
wire mux_o_1985;
wire mux_o_1986;
wire mux_o_1987;
wire mux_o_1988;
wire mux_o_1989;
wire mux_o_1990;
wire mux_o_1991;
wire mux_o_1992;
wire mux_o_1993;
wire mux_o_1994;
wire mux_o_1995;
wire mux_o_1996;
wire mux_o_1997;
wire mux_o_1998;
wire mux_o_1999;
wire mux_o_2000;
wire mux_o_2001;
wire mux_o_2002;
wire mux_o_2003;
wire mux_o_2004;
wire mux_o_2005;
wire mux_o_2006;
wire mux_o_2007;
wire mux_o_2008;
wire mux_o_2009;
wire mux_o_2010;
wire mux_o_2011;
wire mux_o_2012;
wire mux_o_2013;
wire mux_o_2014;
wire mux_o_2015;
wire mux_o_2016;
wire mux_o_2017;
wire mux_o_2018;
wire mux_o_2019;
wire mux_o_2020;
wire mux_o_2021;
wire mux_o_2022;
wire mux_o_2023;
wire mux_o_2024;
wire mux_o_2025;
wire mux_o_2026;
wire mux_o_2027;
wire mux_o_2028;
wire mux_o_2029;
wire mux_o_2030;
wire mux_o_2032;
wire mux_o_2033;
wire mux_o_2034;
wire mux_o_2035;
wire mux_o_2036;
wire mux_o_2037;
wire mux_o_2038;
wire mux_o_2039;
wire mux_o_2040;
wire mux_o_2041;
wire mux_o_2042;
wire mux_o_2043;
wire mux_o_2044;
wire mux_o_2045;
wire mux_o_2046;
wire mux_o_2047;
wire mux_o_2048;
wire mux_o_2049;
wire mux_o_2050;
wire mux_o_2051;
wire mux_o_2052;
wire mux_o_2053;
wire mux_o_2054;
wire mux_o_2055;
wire mux_o_2056;
wire mux_o_2057;
wire mux_o_2058;
wire mux_o_2059;
wire mux_o_2060;
wire mux_o_2061;
wire mux_o_2062;
wire mux_o_2063;
wire mux_o_2064;
wire mux_o_2065;
wire mux_o_2066;
wire mux_o_2067;
wire mux_o_2068;
wire mux_o_2069;
wire mux_o_2070;
wire mux_o_2071;
wire mux_o_2072;
wire mux_o_2073;
wire mux_o_2074;
wire mux_o_2075;
wire mux_o_2076;
wire mux_o_2077;
wire mux_o_2078;
wire mux_o_2079;
wire mux_o_2080;
wire mux_o_2081;
wire mux_o_2082;
wire mux_o_2083;
wire mux_o_2084;
wire mux_o_2085;
wire mux_o_2086;
wire mux_o_2087;
wire mux_o_2088;
wire mux_o_2089;
wire mux_o_2090;
wire mux_o_2091;
wire mux_o_2092;
wire mux_o_2093;
wire mux_o_2094;
wire mux_o_2095;
wire mux_o_2096;
wire mux_o_2097;
wire mux_o_2098;
wire mux_o_2099;
wire mux_o_2100;
wire mux_o_2101;
wire mux_o_2102;
wire mux_o_2103;
wire mux_o_2104;
wire mux_o_2105;
wire mux_o_2106;
wire mux_o_2107;
wire mux_o_2108;
wire mux_o_2109;
wire mux_o_2110;
wire mux_o_2111;
wire mux_o_2112;
wire mux_o_2113;
wire mux_o_2114;
wire mux_o_2115;
wire mux_o_2116;
wire mux_o_2117;
wire mux_o_2118;
wire mux_o_2119;
wire mux_o_2120;
wire mux_o_2121;
wire mux_o_2122;
wire mux_o_2123;
wire mux_o_2124;
wire mux_o_2125;
wire mux_o_2126;
wire mux_o_2127;
wire mux_o_2128;
wire mux_o_2129;
wire mux_o_2130;
wire mux_o_2131;
wire mux_o_2132;
wire mux_o_2133;
wire mux_o_2134;
wire mux_o_2135;
wire mux_o_2136;
wire mux_o_2137;
wire mux_o_2138;
wire mux_o_2139;
wire mux_o_2140;
wire mux_o_2141;
wire mux_o_2142;
wire mux_o_2143;
wire mux_o_2144;
wire mux_o_2145;
wire mux_o_2146;
wire mux_o_2147;
wire mux_o_2148;
wire mux_o_2149;
wire mux_o_2150;
wire mux_o_2151;
wire mux_o_2152;
wire mux_o_2153;
wire mux_o_2154;
wire mux_o_2155;
wire mux_o_2156;
wire mux_o_2157;
wire mux_o_2159;
wire mux_o_2160;
wire mux_o_2161;
wire mux_o_2162;
wire mux_o_2163;
wire mux_o_2164;
wire mux_o_2165;
wire mux_o_2166;
wire mux_o_2167;
wire mux_o_2168;
wire mux_o_2169;
wire mux_o_2170;
wire mux_o_2171;
wire mux_o_2172;
wire mux_o_2173;
wire mux_o_2174;
wire mux_o_2175;
wire mux_o_2176;
wire mux_o_2177;
wire mux_o_2178;
wire mux_o_2179;
wire mux_o_2180;
wire mux_o_2181;
wire mux_o_2182;
wire mux_o_2183;
wire mux_o_2184;
wire mux_o_2185;
wire mux_o_2186;
wire mux_o_2187;
wire mux_o_2188;
wire mux_o_2189;
wire mux_o_2190;
wire mux_o_2191;
wire mux_o_2192;
wire mux_o_2193;
wire mux_o_2194;
wire mux_o_2195;
wire mux_o_2196;
wire mux_o_2197;
wire mux_o_2198;
wire mux_o_2199;
wire mux_o_2200;
wire mux_o_2201;
wire mux_o_2202;
wire mux_o_2203;
wire mux_o_2204;
wire mux_o_2205;
wire mux_o_2206;
wire mux_o_2207;
wire mux_o_2208;
wire mux_o_2209;
wire mux_o_2210;
wire mux_o_2211;
wire mux_o_2212;
wire mux_o_2213;
wire mux_o_2214;
wire mux_o_2215;
wire mux_o_2216;
wire mux_o_2217;
wire mux_o_2218;
wire mux_o_2219;
wire mux_o_2220;
wire mux_o_2221;
wire mux_o_2222;
wire mux_o_2223;
wire mux_o_2224;
wire mux_o_2225;
wire mux_o_2226;
wire mux_o_2227;
wire mux_o_2228;
wire mux_o_2229;
wire mux_o_2230;
wire mux_o_2231;
wire mux_o_2232;
wire mux_o_2233;
wire mux_o_2234;
wire mux_o_2235;
wire mux_o_2236;
wire mux_o_2237;
wire mux_o_2238;
wire mux_o_2239;
wire mux_o_2240;
wire mux_o_2241;
wire mux_o_2242;
wire mux_o_2243;
wire mux_o_2244;
wire mux_o_2245;
wire mux_o_2246;
wire mux_o_2247;
wire mux_o_2248;
wire mux_o_2249;
wire mux_o_2250;
wire mux_o_2251;
wire mux_o_2252;
wire mux_o_2253;
wire mux_o_2254;
wire mux_o_2255;
wire mux_o_2256;
wire mux_o_2257;
wire mux_o_2258;
wire mux_o_2259;
wire mux_o_2260;
wire mux_o_2261;
wire mux_o_2262;
wire mux_o_2263;
wire mux_o_2264;
wire mux_o_2265;
wire mux_o_2266;
wire mux_o_2267;
wire mux_o_2268;
wire mux_o_2269;
wire mux_o_2270;
wire mux_o_2271;
wire mux_o_2272;
wire mux_o_2273;
wire mux_o_2274;
wire mux_o_2275;
wire mux_o_2276;
wire mux_o_2277;
wire mux_o_2278;
wire mux_o_2279;
wire mux_o_2280;
wire mux_o_2281;
wire mux_o_2282;
wire mux_o_2283;
wire mux_o_2284;
wire mux_o_2286;
wire mux_o_2287;
wire mux_o_2288;
wire mux_o_2289;
wire mux_o_2290;
wire mux_o_2291;
wire mux_o_2292;
wire mux_o_2293;
wire mux_o_2294;
wire mux_o_2295;
wire mux_o_2296;
wire mux_o_2297;
wire mux_o_2298;
wire mux_o_2299;
wire mux_o_2300;
wire mux_o_2301;
wire mux_o_2302;
wire mux_o_2303;
wire mux_o_2304;
wire mux_o_2305;
wire mux_o_2306;
wire mux_o_2307;
wire mux_o_2308;
wire mux_o_2309;
wire mux_o_2310;
wire mux_o_2311;
wire mux_o_2312;
wire mux_o_2313;
wire mux_o_2314;
wire mux_o_2315;
wire mux_o_2316;
wire mux_o_2317;
wire mux_o_2318;
wire mux_o_2319;
wire mux_o_2320;
wire mux_o_2321;
wire mux_o_2322;
wire mux_o_2323;
wire mux_o_2324;
wire mux_o_2325;
wire mux_o_2326;
wire mux_o_2327;
wire mux_o_2328;
wire mux_o_2329;
wire mux_o_2330;
wire mux_o_2331;
wire mux_o_2332;
wire mux_o_2333;
wire mux_o_2334;
wire mux_o_2335;
wire mux_o_2336;
wire mux_o_2337;
wire mux_o_2338;
wire mux_o_2339;
wire mux_o_2340;
wire mux_o_2341;
wire mux_o_2342;
wire mux_o_2343;
wire mux_o_2344;
wire mux_o_2345;
wire mux_o_2346;
wire mux_o_2347;
wire mux_o_2348;
wire mux_o_2349;
wire mux_o_2350;
wire mux_o_2351;
wire mux_o_2352;
wire mux_o_2353;
wire mux_o_2354;
wire mux_o_2355;
wire mux_o_2356;
wire mux_o_2357;
wire mux_o_2358;
wire mux_o_2359;
wire mux_o_2360;
wire mux_o_2361;
wire mux_o_2362;
wire mux_o_2363;
wire mux_o_2364;
wire mux_o_2365;
wire mux_o_2366;
wire mux_o_2367;
wire mux_o_2368;
wire mux_o_2369;
wire mux_o_2370;
wire mux_o_2371;
wire mux_o_2372;
wire mux_o_2373;
wire mux_o_2374;
wire mux_o_2375;
wire mux_o_2376;
wire mux_o_2377;
wire mux_o_2378;
wire mux_o_2379;
wire mux_o_2380;
wire mux_o_2381;
wire mux_o_2382;
wire mux_o_2383;
wire mux_o_2384;
wire mux_o_2385;
wire mux_o_2386;
wire mux_o_2387;
wire mux_o_2388;
wire mux_o_2389;
wire mux_o_2390;
wire mux_o_2391;
wire mux_o_2392;
wire mux_o_2393;
wire mux_o_2394;
wire mux_o_2395;
wire mux_o_2396;
wire mux_o_2397;
wire mux_o_2398;
wire mux_o_2399;
wire mux_o_2400;
wire mux_o_2401;
wire mux_o_2402;
wire mux_o_2403;
wire mux_o_2404;
wire mux_o_2405;
wire mux_o_2406;
wire mux_o_2407;
wire mux_o_2408;
wire mux_o_2409;
wire mux_o_2410;
wire mux_o_2411;
wire mux_o_2413;
wire mux_o_2414;
wire mux_o_2415;
wire mux_o_2416;
wire mux_o_2417;
wire mux_o_2418;
wire mux_o_2419;
wire mux_o_2420;
wire mux_o_2421;
wire mux_o_2422;
wire mux_o_2423;
wire mux_o_2424;
wire mux_o_2425;
wire mux_o_2426;
wire mux_o_2427;
wire mux_o_2428;
wire mux_o_2429;
wire mux_o_2430;
wire mux_o_2431;
wire mux_o_2432;
wire mux_o_2433;
wire mux_o_2434;
wire mux_o_2435;
wire mux_o_2436;
wire mux_o_2437;
wire mux_o_2438;
wire mux_o_2439;
wire mux_o_2440;
wire mux_o_2441;
wire mux_o_2442;
wire mux_o_2443;
wire mux_o_2444;
wire mux_o_2445;
wire mux_o_2446;
wire mux_o_2447;
wire mux_o_2448;
wire mux_o_2449;
wire mux_o_2450;
wire mux_o_2451;
wire mux_o_2452;
wire mux_o_2453;
wire mux_o_2454;
wire mux_o_2455;
wire mux_o_2456;
wire mux_o_2457;
wire mux_o_2458;
wire mux_o_2459;
wire mux_o_2460;
wire mux_o_2461;
wire mux_o_2462;
wire mux_o_2463;
wire mux_o_2464;
wire mux_o_2465;
wire mux_o_2466;
wire mux_o_2467;
wire mux_o_2468;
wire mux_o_2469;
wire mux_o_2470;
wire mux_o_2471;
wire mux_o_2472;
wire mux_o_2473;
wire mux_o_2474;
wire mux_o_2475;
wire mux_o_2476;
wire mux_o_2477;
wire mux_o_2478;
wire mux_o_2479;
wire mux_o_2480;
wire mux_o_2481;
wire mux_o_2482;
wire mux_o_2483;
wire mux_o_2484;
wire mux_o_2485;
wire mux_o_2486;
wire mux_o_2487;
wire mux_o_2488;
wire mux_o_2489;
wire mux_o_2490;
wire mux_o_2491;
wire mux_o_2492;
wire mux_o_2493;
wire mux_o_2494;
wire mux_o_2495;
wire mux_o_2496;
wire mux_o_2497;
wire mux_o_2498;
wire mux_o_2499;
wire mux_o_2500;
wire mux_o_2501;
wire mux_o_2502;
wire mux_o_2503;
wire mux_o_2504;
wire mux_o_2505;
wire mux_o_2506;
wire mux_o_2507;
wire mux_o_2508;
wire mux_o_2509;
wire mux_o_2510;
wire mux_o_2511;
wire mux_o_2512;
wire mux_o_2513;
wire mux_o_2514;
wire mux_o_2515;
wire mux_o_2516;
wire mux_o_2517;
wire mux_o_2518;
wire mux_o_2519;
wire mux_o_2520;
wire mux_o_2521;
wire mux_o_2522;
wire mux_o_2523;
wire mux_o_2524;
wire mux_o_2525;
wire mux_o_2526;
wire mux_o_2527;
wire mux_o_2528;
wire mux_o_2529;
wire mux_o_2530;
wire mux_o_2531;
wire mux_o_2532;
wire mux_o_2533;
wire mux_o_2534;
wire mux_o_2535;
wire mux_o_2536;
wire mux_o_2537;
wire mux_o_2538;
wire mux_o_2540;
wire mux_o_2541;
wire mux_o_2542;
wire mux_o_2543;
wire mux_o_2544;
wire mux_o_2545;
wire mux_o_2546;
wire mux_o_2547;
wire mux_o_2548;
wire mux_o_2549;
wire mux_o_2550;
wire mux_o_2551;
wire mux_o_2552;
wire mux_o_2553;
wire mux_o_2554;
wire mux_o_2555;
wire mux_o_2556;
wire mux_o_2557;
wire mux_o_2558;
wire mux_o_2559;
wire mux_o_2560;
wire mux_o_2561;
wire mux_o_2562;
wire mux_o_2563;
wire mux_o_2564;
wire mux_o_2565;
wire mux_o_2566;
wire mux_o_2567;
wire mux_o_2568;
wire mux_o_2569;
wire mux_o_2570;
wire mux_o_2571;
wire mux_o_2572;
wire mux_o_2573;
wire mux_o_2574;
wire mux_o_2575;
wire mux_o_2576;
wire mux_o_2577;
wire mux_o_2578;
wire mux_o_2579;
wire mux_o_2580;
wire mux_o_2581;
wire mux_o_2582;
wire mux_o_2583;
wire mux_o_2584;
wire mux_o_2585;
wire mux_o_2586;
wire mux_o_2587;
wire mux_o_2588;
wire mux_o_2589;
wire mux_o_2590;
wire mux_o_2591;
wire mux_o_2592;
wire mux_o_2593;
wire mux_o_2594;
wire mux_o_2595;
wire mux_o_2596;
wire mux_o_2597;
wire mux_o_2598;
wire mux_o_2599;
wire mux_o_2600;
wire mux_o_2601;
wire mux_o_2602;
wire mux_o_2603;
wire mux_o_2604;
wire mux_o_2605;
wire mux_o_2606;
wire mux_o_2607;
wire mux_o_2608;
wire mux_o_2609;
wire mux_o_2610;
wire mux_o_2611;
wire mux_o_2612;
wire mux_o_2613;
wire mux_o_2614;
wire mux_o_2615;
wire mux_o_2616;
wire mux_o_2617;
wire mux_o_2618;
wire mux_o_2619;
wire mux_o_2620;
wire mux_o_2621;
wire mux_o_2622;
wire mux_o_2623;
wire mux_o_2624;
wire mux_o_2625;
wire mux_o_2626;
wire mux_o_2627;
wire mux_o_2628;
wire mux_o_2629;
wire mux_o_2630;
wire mux_o_2631;
wire mux_o_2632;
wire mux_o_2633;
wire mux_o_2634;
wire mux_o_2635;
wire mux_o_2636;
wire mux_o_2637;
wire mux_o_2638;
wire mux_o_2639;
wire mux_o_2640;
wire mux_o_2641;
wire mux_o_2642;
wire mux_o_2643;
wire mux_o_2644;
wire mux_o_2645;
wire mux_o_2646;
wire mux_o_2647;
wire mux_o_2648;
wire mux_o_2649;
wire mux_o_2650;
wire mux_o_2651;
wire mux_o_2652;
wire mux_o_2653;
wire mux_o_2654;
wire mux_o_2655;
wire mux_o_2656;
wire mux_o_2657;
wire mux_o_2658;
wire mux_o_2659;
wire mux_o_2660;
wire mux_o_2661;
wire mux_o_2662;
wire mux_o_2663;
wire mux_o_2664;
wire mux_o_2665;
wire mux_o_2667;
wire mux_o_2668;
wire mux_o_2669;
wire mux_o_2670;
wire mux_o_2671;
wire mux_o_2672;
wire mux_o_2673;
wire mux_o_2674;
wire mux_o_2675;
wire mux_o_2676;
wire mux_o_2677;
wire mux_o_2678;
wire mux_o_2679;
wire mux_o_2680;
wire mux_o_2681;
wire mux_o_2682;
wire mux_o_2683;
wire mux_o_2684;
wire mux_o_2685;
wire mux_o_2686;
wire mux_o_2687;
wire mux_o_2688;
wire mux_o_2689;
wire mux_o_2690;
wire mux_o_2691;
wire mux_o_2692;
wire mux_o_2693;
wire mux_o_2694;
wire mux_o_2695;
wire mux_o_2696;
wire mux_o_2697;
wire mux_o_2698;
wire mux_o_2699;
wire mux_o_2700;
wire mux_o_2701;
wire mux_o_2702;
wire mux_o_2703;
wire mux_o_2704;
wire mux_o_2705;
wire mux_o_2706;
wire mux_o_2707;
wire mux_o_2708;
wire mux_o_2709;
wire mux_o_2710;
wire mux_o_2711;
wire mux_o_2712;
wire mux_o_2713;
wire mux_o_2714;
wire mux_o_2715;
wire mux_o_2716;
wire mux_o_2717;
wire mux_o_2718;
wire mux_o_2719;
wire mux_o_2720;
wire mux_o_2721;
wire mux_o_2722;
wire mux_o_2723;
wire mux_o_2724;
wire mux_o_2725;
wire mux_o_2726;
wire mux_o_2727;
wire mux_o_2728;
wire mux_o_2729;
wire mux_o_2730;
wire mux_o_2731;
wire mux_o_2732;
wire mux_o_2733;
wire mux_o_2734;
wire mux_o_2735;
wire mux_o_2736;
wire mux_o_2737;
wire mux_o_2738;
wire mux_o_2739;
wire mux_o_2740;
wire mux_o_2741;
wire mux_o_2742;
wire mux_o_2743;
wire mux_o_2744;
wire mux_o_2745;
wire mux_o_2746;
wire mux_o_2747;
wire mux_o_2748;
wire mux_o_2749;
wire mux_o_2750;
wire mux_o_2751;
wire mux_o_2752;
wire mux_o_2753;
wire mux_o_2754;
wire mux_o_2755;
wire mux_o_2756;
wire mux_o_2757;
wire mux_o_2758;
wire mux_o_2759;
wire mux_o_2760;
wire mux_o_2761;
wire mux_o_2762;
wire mux_o_2763;
wire mux_o_2764;
wire mux_o_2765;
wire mux_o_2766;
wire mux_o_2767;
wire mux_o_2768;
wire mux_o_2769;
wire mux_o_2770;
wire mux_o_2771;
wire mux_o_2772;
wire mux_o_2773;
wire mux_o_2774;
wire mux_o_2775;
wire mux_o_2776;
wire mux_o_2777;
wire mux_o_2778;
wire mux_o_2779;
wire mux_o_2780;
wire mux_o_2781;
wire mux_o_2782;
wire mux_o_2783;
wire mux_o_2784;
wire mux_o_2785;
wire mux_o_2786;
wire mux_o_2787;
wire mux_o_2788;
wire mux_o_2789;
wire mux_o_2790;
wire mux_o_2791;
wire mux_o_2792;
wire mux_o_2794;
wire mux_o_2795;
wire mux_o_2796;
wire mux_o_2797;
wire mux_o_2798;
wire mux_o_2799;
wire mux_o_2800;
wire mux_o_2801;
wire mux_o_2802;
wire mux_o_2803;
wire mux_o_2804;
wire mux_o_2805;
wire mux_o_2806;
wire mux_o_2807;
wire mux_o_2808;
wire mux_o_2809;
wire mux_o_2810;
wire mux_o_2811;
wire mux_o_2812;
wire mux_o_2813;
wire mux_o_2814;
wire mux_o_2815;
wire mux_o_2816;
wire mux_o_2817;
wire mux_o_2818;
wire mux_o_2819;
wire mux_o_2820;
wire mux_o_2821;
wire mux_o_2822;
wire mux_o_2823;
wire mux_o_2824;
wire mux_o_2825;
wire mux_o_2826;
wire mux_o_2827;
wire mux_o_2828;
wire mux_o_2829;
wire mux_o_2830;
wire mux_o_2831;
wire mux_o_2832;
wire mux_o_2833;
wire mux_o_2834;
wire mux_o_2835;
wire mux_o_2836;
wire mux_o_2837;
wire mux_o_2838;
wire mux_o_2839;
wire mux_o_2840;
wire mux_o_2841;
wire mux_o_2842;
wire mux_o_2843;
wire mux_o_2844;
wire mux_o_2845;
wire mux_o_2846;
wire mux_o_2847;
wire mux_o_2848;
wire mux_o_2849;
wire mux_o_2850;
wire mux_o_2851;
wire mux_o_2852;
wire mux_o_2853;
wire mux_o_2854;
wire mux_o_2855;
wire mux_o_2856;
wire mux_o_2857;
wire mux_o_2858;
wire mux_o_2859;
wire mux_o_2860;
wire mux_o_2861;
wire mux_o_2862;
wire mux_o_2863;
wire mux_o_2864;
wire mux_o_2865;
wire mux_o_2866;
wire mux_o_2867;
wire mux_o_2868;
wire mux_o_2869;
wire mux_o_2870;
wire mux_o_2871;
wire mux_o_2872;
wire mux_o_2873;
wire mux_o_2874;
wire mux_o_2875;
wire mux_o_2876;
wire mux_o_2877;
wire mux_o_2878;
wire mux_o_2879;
wire mux_o_2880;
wire mux_o_2881;
wire mux_o_2882;
wire mux_o_2883;
wire mux_o_2884;
wire mux_o_2885;
wire mux_o_2886;
wire mux_o_2887;
wire mux_o_2888;
wire mux_o_2889;
wire mux_o_2890;
wire mux_o_2891;
wire mux_o_2892;
wire mux_o_2893;
wire mux_o_2894;
wire mux_o_2895;
wire mux_o_2896;
wire mux_o_2897;
wire mux_o_2898;
wire mux_o_2899;
wire mux_o_2900;
wire mux_o_2901;
wire mux_o_2902;
wire mux_o_2903;
wire mux_o_2904;
wire mux_o_2905;
wire mux_o_2906;
wire mux_o_2907;
wire mux_o_2908;
wire mux_o_2909;
wire mux_o_2910;
wire mux_o_2911;
wire mux_o_2912;
wire mux_o_2913;
wire mux_o_2914;
wire mux_o_2915;
wire mux_o_2916;
wire mux_o_2917;
wire mux_o_2918;
wire mux_o_2919;
wire mux_o_2921;
wire mux_o_2922;
wire mux_o_2923;
wire mux_o_2924;
wire mux_o_2925;
wire mux_o_2926;
wire mux_o_2927;
wire mux_o_2928;
wire mux_o_2929;
wire mux_o_2930;
wire mux_o_2931;
wire mux_o_2932;
wire mux_o_2933;
wire mux_o_2934;
wire mux_o_2935;
wire mux_o_2936;
wire mux_o_2937;
wire mux_o_2938;
wire mux_o_2939;
wire mux_o_2940;
wire mux_o_2941;
wire mux_o_2942;
wire mux_o_2943;
wire mux_o_2944;
wire mux_o_2945;
wire mux_o_2946;
wire mux_o_2947;
wire mux_o_2948;
wire mux_o_2949;
wire mux_o_2950;
wire mux_o_2951;
wire mux_o_2952;
wire mux_o_2953;
wire mux_o_2954;
wire mux_o_2955;
wire mux_o_2956;
wire mux_o_2957;
wire mux_o_2958;
wire mux_o_2959;
wire mux_o_2960;
wire mux_o_2961;
wire mux_o_2962;
wire mux_o_2963;
wire mux_o_2964;
wire mux_o_2965;
wire mux_o_2966;
wire mux_o_2967;
wire mux_o_2968;
wire mux_o_2969;
wire mux_o_2970;
wire mux_o_2971;
wire mux_o_2972;
wire mux_o_2973;
wire mux_o_2974;
wire mux_o_2975;
wire mux_o_2976;
wire mux_o_2977;
wire mux_o_2978;
wire mux_o_2979;
wire mux_o_2980;
wire mux_o_2981;
wire mux_o_2982;
wire mux_o_2983;
wire mux_o_2984;
wire mux_o_2985;
wire mux_o_2986;
wire mux_o_2987;
wire mux_o_2988;
wire mux_o_2989;
wire mux_o_2990;
wire mux_o_2991;
wire mux_o_2992;
wire mux_o_2993;
wire mux_o_2994;
wire mux_o_2995;
wire mux_o_2996;
wire mux_o_2997;
wire mux_o_2998;
wire mux_o_2999;
wire mux_o_3000;
wire mux_o_3001;
wire mux_o_3002;
wire mux_o_3003;
wire mux_o_3004;
wire mux_o_3005;
wire mux_o_3006;
wire mux_o_3007;
wire mux_o_3008;
wire mux_o_3009;
wire mux_o_3010;
wire mux_o_3011;
wire mux_o_3012;
wire mux_o_3013;
wire mux_o_3014;
wire mux_o_3015;
wire mux_o_3016;
wire mux_o_3017;
wire mux_o_3018;
wire mux_o_3019;
wire mux_o_3020;
wire mux_o_3021;
wire mux_o_3022;
wire mux_o_3023;
wire mux_o_3024;
wire mux_o_3025;
wire mux_o_3026;
wire mux_o_3027;
wire mux_o_3028;
wire mux_o_3029;
wire mux_o_3030;
wire mux_o_3031;
wire mux_o_3032;
wire mux_o_3033;
wire mux_o_3034;
wire mux_o_3035;
wire mux_o_3036;
wire mux_o_3037;
wire mux_o_3038;
wire mux_o_3039;
wire mux_o_3040;
wire mux_o_3041;
wire mux_o_3042;
wire mux_o_3043;
wire mux_o_3044;
wire mux_o_3045;
wire mux_o_3046;
wire mux_o_3048;
wire mux_o_3049;
wire mux_o_3050;
wire mux_o_3051;
wire mux_o_3052;
wire mux_o_3053;
wire mux_o_3054;
wire mux_o_3055;
wire mux_o_3056;
wire mux_o_3057;
wire mux_o_3058;
wire mux_o_3059;
wire mux_o_3060;
wire mux_o_3061;
wire mux_o_3062;
wire mux_o_3063;
wire mux_o_3064;
wire mux_o_3065;
wire mux_o_3066;
wire mux_o_3067;
wire mux_o_3068;
wire mux_o_3069;
wire mux_o_3070;
wire mux_o_3071;
wire mux_o_3072;
wire mux_o_3073;
wire mux_o_3074;
wire mux_o_3075;
wire mux_o_3076;
wire mux_o_3077;
wire mux_o_3078;
wire mux_o_3079;
wire mux_o_3080;
wire mux_o_3081;
wire mux_o_3082;
wire mux_o_3083;
wire mux_o_3084;
wire mux_o_3085;
wire mux_o_3086;
wire mux_o_3087;
wire mux_o_3088;
wire mux_o_3089;
wire mux_o_3090;
wire mux_o_3091;
wire mux_o_3092;
wire mux_o_3093;
wire mux_o_3094;
wire mux_o_3095;
wire mux_o_3096;
wire mux_o_3097;
wire mux_o_3098;
wire mux_o_3099;
wire mux_o_3100;
wire mux_o_3101;
wire mux_o_3102;
wire mux_o_3103;
wire mux_o_3104;
wire mux_o_3105;
wire mux_o_3106;
wire mux_o_3107;
wire mux_o_3108;
wire mux_o_3109;
wire mux_o_3110;
wire mux_o_3111;
wire mux_o_3112;
wire mux_o_3113;
wire mux_o_3114;
wire mux_o_3115;
wire mux_o_3116;
wire mux_o_3117;
wire mux_o_3118;
wire mux_o_3119;
wire mux_o_3120;
wire mux_o_3121;
wire mux_o_3122;
wire mux_o_3123;
wire mux_o_3124;
wire mux_o_3125;
wire mux_o_3126;
wire mux_o_3127;
wire mux_o_3128;
wire mux_o_3129;
wire mux_o_3130;
wire mux_o_3131;
wire mux_o_3132;
wire mux_o_3133;
wire mux_o_3134;
wire mux_o_3135;
wire mux_o_3136;
wire mux_o_3137;
wire mux_o_3138;
wire mux_o_3139;
wire mux_o_3140;
wire mux_o_3141;
wire mux_o_3142;
wire mux_o_3143;
wire mux_o_3144;
wire mux_o_3145;
wire mux_o_3146;
wire mux_o_3147;
wire mux_o_3148;
wire mux_o_3149;
wire mux_o_3150;
wire mux_o_3151;
wire mux_o_3152;
wire mux_o_3153;
wire mux_o_3154;
wire mux_o_3155;
wire mux_o_3156;
wire mux_o_3157;
wire mux_o_3158;
wire mux_o_3159;
wire mux_o_3160;
wire mux_o_3161;
wire mux_o_3162;
wire mux_o_3163;
wire mux_o_3164;
wire mux_o_3165;
wire mux_o_3166;
wire mux_o_3167;
wire mux_o_3168;
wire mux_o_3169;
wire mux_o_3170;
wire mux_o_3171;
wire mux_o_3172;
wire mux_o_3173;
wire mux_o_3175;
wire mux_o_3176;
wire mux_o_3177;
wire mux_o_3178;
wire mux_o_3179;
wire mux_o_3180;
wire mux_o_3181;
wire mux_o_3182;
wire mux_o_3183;
wire mux_o_3184;
wire mux_o_3185;
wire mux_o_3186;
wire mux_o_3187;
wire mux_o_3188;
wire mux_o_3189;
wire mux_o_3190;
wire mux_o_3191;
wire mux_o_3192;
wire mux_o_3193;
wire mux_o_3194;
wire mux_o_3195;
wire mux_o_3196;
wire mux_o_3197;
wire mux_o_3198;
wire mux_o_3199;
wire mux_o_3200;
wire mux_o_3201;
wire mux_o_3202;
wire mux_o_3203;
wire mux_o_3204;
wire mux_o_3205;
wire mux_o_3206;
wire mux_o_3207;
wire mux_o_3208;
wire mux_o_3209;
wire mux_o_3210;
wire mux_o_3211;
wire mux_o_3212;
wire mux_o_3213;
wire mux_o_3214;
wire mux_o_3215;
wire mux_o_3216;
wire mux_o_3217;
wire mux_o_3218;
wire mux_o_3219;
wire mux_o_3220;
wire mux_o_3221;
wire mux_o_3222;
wire mux_o_3223;
wire mux_o_3224;
wire mux_o_3225;
wire mux_o_3226;
wire mux_o_3227;
wire mux_o_3228;
wire mux_o_3229;
wire mux_o_3230;
wire mux_o_3231;
wire mux_o_3232;
wire mux_o_3233;
wire mux_o_3234;
wire mux_o_3235;
wire mux_o_3236;
wire mux_o_3237;
wire mux_o_3238;
wire mux_o_3239;
wire mux_o_3240;
wire mux_o_3241;
wire mux_o_3242;
wire mux_o_3243;
wire mux_o_3244;
wire mux_o_3245;
wire mux_o_3246;
wire mux_o_3247;
wire mux_o_3248;
wire mux_o_3249;
wire mux_o_3250;
wire mux_o_3251;
wire mux_o_3252;
wire mux_o_3253;
wire mux_o_3254;
wire mux_o_3255;
wire mux_o_3256;
wire mux_o_3257;
wire mux_o_3258;
wire mux_o_3259;
wire mux_o_3260;
wire mux_o_3261;
wire mux_o_3262;
wire mux_o_3263;
wire mux_o_3264;
wire mux_o_3265;
wire mux_o_3266;
wire mux_o_3267;
wire mux_o_3268;
wire mux_o_3269;
wire mux_o_3270;
wire mux_o_3271;
wire mux_o_3272;
wire mux_o_3273;
wire mux_o_3274;
wire mux_o_3275;
wire mux_o_3276;
wire mux_o_3277;
wire mux_o_3278;
wire mux_o_3279;
wire mux_o_3280;
wire mux_o_3281;
wire mux_o_3282;
wire mux_o_3283;
wire mux_o_3284;
wire mux_o_3285;
wire mux_o_3286;
wire mux_o_3287;
wire mux_o_3288;
wire mux_o_3289;
wire mux_o_3290;
wire mux_o_3291;
wire mux_o_3292;
wire mux_o_3293;
wire mux_o_3294;
wire mux_o_3295;
wire mux_o_3296;
wire mux_o_3297;
wire mux_o_3298;
wire mux_o_3299;
wire mux_o_3300;
wire mux_o_3302;
wire mux_o_3303;
wire mux_o_3304;
wire mux_o_3305;
wire mux_o_3306;
wire mux_o_3307;
wire mux_o_3308;
wire mux_o_3309;
wire mux_o_3310;
wire mux_o_3311;
wire mux_o_3312;
wire mux_o_3313;
wire mux_o_3314;
wire mux_o_3315;
wire mux_o_3316;
wire mux_o_3317;
wire mux_o_3318;
wire mux_o_3319;
wire mux_o_3320;
wire mux_o_3321;
wire mux_o_3322;
wire mux_o_3323;
wire mux_o_3324;
wire mux_o_3325;
wire mux_o_3326;
wire mux_o_3327;
wire mux_o_3328;
wire mux_o_3329;
wire mux_o_3330;
wire mux_o_3331;
wire mux_o_3332;
wire mux_o_3333;
wire mux_o_3334;
wire mux_o_3335;
wire mux_o_3336;
wire mux_o_3337;
wire mux_o_3338;
wire mux_o_3339;
wire mux_o_3340;
wire mux_o_3341;
wire mux_o_3342;
wire mux_o_3343;
wire mux_o_3344;
wire mux_o_3345;
wire mux_o_3346;
wire mux_o_3347;
wire mux_o_3348;
wire mux_o_3349;
wire mux_o_3350;
wire mux_o_3351;
wire mux_o_3352;
wire mux_o_3353;
wire mux_o_3354;
wire mux_o_3355;
wire mux_o_3356;
wire mux_o_3357;
wire mux_o_3358;
wire mux_o_3359;
wire mux_o_3360;
wire mux_o_3361;
wire mux_o_3362;
wire mux_o_3363;
wire mux_o_3364;
wire mux_o_3365;
wire mux_o_3366;
wire mux_o_3367;
wire mux_o_3368;
wire mux_o_3369;
wire mux_o_3370;
wire mux_o_3371;
wire mux_o_3372;
wire mux_o_3373;
wire mux_o_3374;
wire mux_o_3375;
wire mux_o_3376;
wire mux_o_3377;
wire mux_o_3378;
wire mux_o_3379;
wire mux_o_3380;
wire mux_o_3381;
wire mux_o_3382;
wire mux_o_3383;
wire mux_o_3384;
wire mux_o_3385;
wire mux_o_3386;
wire mux_o_3387;
wire mux_o_3388;
wire mux_o_3389;
wire mux_o_3390;
wire mux_o_3391;
wire mux_o_3392;
wire mux_o_3393;
wire mux_o_3394;
wire mux_o_3395;
wire mux_o_3396;
wire mux_o_3397;
wire mux_o_3398;
wire mux_o_3399;
wire mux_o_3400;
wire mux_o_3401;
wire mux_o_3402;
wire mux_o_3403;
wire mux_o_3404;
wire mux_o_3405;
wire mux_o_3406;
wire mux_o_3407;
wire mux_o_3408;
wire mux_o_3409;
wire mux_o_3410;
wire mux_o_3411;
wire mux_o_3412;
wire mux_o_3413;
wire mux_o_3414;
wire mux_o_3415;
wire mux_o_3416;
wire mux_o_3417;
wire mux_o_3418;
wire mux_o_3419;
wire mux_o_3420;
wire mux_o_3421;
wire mux_o_3422;
wire mux_o_3423;
wire mux_o_3424;
wire mux_o_3425;
wire mux_o_3426;
wire mux_o_3427;
wire mux_o_3429;
wire mux_o_3430;
wire mux_o_3431;
wire mux_o_3432;
wire mux_o_3433;
wire mux_o_3434;
wire mux_o_3435;
wire mux_o_3436;
wire mux_o_3437;
wire mux_o_3438;
wire mux_o_3439;
wire mux_o_3440;
wire mux_o_3441;
wire mux_o_3442;
wire mux_o_3443;
wire mux_o_3444;
wire mux_o_3445;
wire mux_o_3446;
wire mux_o_3447;
wire mux_o_3448;
wire mux_o_3449;
wire mux_o_3450;
wire mux_o_3451;
wire mux_o_3452;
wire mux_o_3453;
wire mux_o_3454;
wire mux_o_3455;
wire mux_o_3456;
wire mux_o_3457;
wire mux_o_3458;
wire mux_o_3459;
wire mux_o_3460;
wire mux_o_3461;
wire mux_o_3462;
wire mux_o_3463;
wire mux_o_3464;
wire mux_o_3465;
wire mux_o_3466;
wire mux_o_3467;
wire mux_o_3468;
wire mux_o_3469;
wire mux_o_3470;
wire mux_o_3471;
wire mux_o_3472;
wire mux_o_3473;
wire mux_o_3474;
wire mux_o_3475;
wire mux_o_3476;
wire mux_o_3477;
wire mux_o_3478;
wire mux_o_3479;
wire mux_o_3480;
wire mux_o_3481;
wire mux_o_3482;
wire mux_o_3483;
wire mux_o_3484;
wire mux_o_3485;
wire mux_o_3486;
wire mux_o_3487;
wire mux_o_3488;
wire mux_o_3489;
wire mux_o_3490;
wire mux_o_3491;
wire mux_o_3492;
wire mux_o_3493;
wire mux_o_3494;
wire mux_o_3495;
wire mux_o_3496;
wire mux_o_3497;
wire mux_o_3498;
wire mux_o_3499;
wire mux_o_3500;
wire mux_o_3501;
wire mux_o_3502;
wire mux_o_3503;
wire mux_o_3504;
wire mux_o_3505;
wire mux_o_3506;
wire mux_o_3507;
wire mux_o_3508;
wire mux_o_3509;
wire mux_o_3510;
wire mux_o_3511;
wire mux_o_3512;
wire mux_o_3513;
wire mux_o_3514;
wire mux_o_3515;
wire mux_o_3516;
wire mux_o_3517;
wire mux_o_3518;
wire mux_o_3519;
wire mux_o_3520;
wire mux_o_3521;
wire mux_o_3522;
wire mux_o_3523;
wire mux_o_3524;
wire mux_o_3525;
wire mux_o_3526;
wire mux_o_3527;
wire mux_o_3528;
wire mux_o_3529;
wire mux_o_3530;
wire mux_o_3531;
wire mux_o_3532;
wire mux_o_3533;
wire mux_o_3534;
wire mux_o_3535;
wire mux_o_3536;
wire mux_o_3537;
wire mux_o_3538;
wire mux_o_3539;
wire mux_o_3540;
wire mux_o_3541;
wire mux_o_3542;
wire mux_o_3543;
wire mux_o_3544;
wire mux_o_3545;
wire mux_o_3546;
wire mux_o_3547;
wire mux_o_3548;
wire mux_o_3549;
wire mux_o_3550;
wire mux_o_3551;
wire mux_o_3552;
wire mux_o_3553;
wire mux_o_3554;
wire mux_o_3556;
wire mux_o_3557;
wire mux_o_3558;
wire mux_o_3559;
wire mux_o_3560;
wire mux_o_3561;
wire mux_o_3562;
wire mux_o_3563;
wire mux_o_3564;
wire mux_o_3565;
wire mux_o_3566;
wire mux_o_3567;
wire mux_o_3568;
wire mux_o_3569;
wire mux_o_3570;
wire mux_o_3571;
wire mux_o_3572;
wire mux_o_3573;
wire mux_o_3574;
wire mux_o_3575;
wire mux_o_3576;
wire mux_o_3577;
wire mux_o_3578;
wire mux_o_3579;
wire mux_o_3580;
wire mux_o_3581;
wire mux_o_3582;
wire mux_o_3583;
wire mux_o_3584;
wire mux_o_3585;
wire mux_o_3586;
wire mux_o_3587;
wire mux_o_3588;
wire mux_o_3589;
wire mux_o_3590;
wire mux_o_3591;
wire mux_o_3592;
wire mux_o_3593;
wire mux_o_3594;
wire mux_o_3595;
wire mux_o_3596;
wire mux_o_3597;
wire mux_o_3598;
wire mux_o_3599;
wire mux_o_3600;
wire mux_o_3601;
wire mux_o_3602;
wire mux_o_3603;
wire mux_o_3604;
wire mux_o_3605;
wire mux_o_3606;
wire mux_o_3607;
wire mux_o_3608;
wire mux_o_3609;
wire mux_o_3610;
wire mux_o_3611;
wire mux_o_3612;
wire mux_o_3613;
wire mux_o_3614;
wire mux_o_3615;
wire mux_o_3616;
wire mux_o_3617;
wire mux_o_3618;
wire mux_o_3619;
wire mux_o_3620;
wire mux_o_3621;
wire mux_o_3622;
wire mux_o_3623;
wire mux_o_3624;
wire mux_o_3625;
wire mux_o_3626;
wire mux_o_3627;
wire mux_o_3628;
wire mux_o_3629;
wire mux_o_3630;
wire mux_o_3631;
wire mux_o_3632;
wire mux_o_3633;
wire mux_o_3634;
wire mux_o_3635;
wire mux_o_3636;
wire mux_o_3637;
wire mux_o_3638;
wire mux_o_3639;
wire mux_o_3640;
wire mux_o_3641;
wire mux_o_3642;
wire mux_o_3643;
wire mux_o_3644;
wire mux_o_3645;
wire mux_o_3646;
wire mux_o_3647;
wire mux_o_3648;
wire mux_o_3649;
wire mux_o_3650;
wire mux_o_3651;
wire mux_o_3652;
wire mux_o_3653;
wire mux_o_3654;
wire mux_o_3655;
wire mux_o_3656;
wire mux_o_3657;
wire mux_o_3658;
wire mux_o_3659;
wire mux_o_3660;
wire mux_o_3661;
wire mux_o_3662;
wire mux_o_3663;
wire mux_o_3664;
wire mux_o_3665;
wire mux_o_3666;
wire mux_o_3667;
wire mux_o_3668;
wire mux_o_3669;
wire mux_o_3670;
wire mux_o_3671;
wire mux_o_3672;
wire mux_o_3673;
wire mux_o_3674;
wire mux_o_3675;
wire mux_o_3676;
wire mux_o_3677;
wire mux_o_3678;
wire mux_o_3679;
wire mux_o_3680;
wire mux_o_3681;
wire mux_o_3683;
wire mux_o_3684;
wire mux_o_3685;
wire mux_o_3686;
wire mux_o_3687;
wire mux_o_3688;
wire mux_o_3689;
wire mux_o_3690;
wire mux_o_3691;
wire mux_o_3692;
wire mux_o_3693;
wire mux_o_3694;
wire mux_o_3695;
wire mux_o_3696;
wire mux_o_3697;
wire mux_o_3698;
wire mux_o_3699;
wire mux_o_3700;
wire mux_o_3701;
wire mux_o_3702;
wire mux_o_3703;
wire mux_o_3704;
wire mux_o_3705;
wire mux_o_3706;
wire mux_o_3707;
wire mux_o_3708;
wire mux_o_3709;
wire mux_o_3710;
wire mux_o_3711;
wire mux_o_3712;
wire mux_o_3713;
wire mux_o_3714;
wire mux_o_3715;
wire mux_o_3716;
wire mux_o_3717;
wire mux_o_3718;
wire mux_o_3719;
wire mux_o_3720;
wire mux_o_3721;
wire mux_o_3722;
wire mux_o_3723;
wire mux_o_3724;
wire mux_o_3725;
wire mux_o_3726;
wire mux_o_3727;
wire mux_o_3728;
wire mux_o_3729;
wire mux_o_3730;
wire mux_o_3731;
wire mux_o_3732;
wire mux_o_3733;
wire mux_o_3734;
wire mux_o_3735;
wire mux_o_3736;
wire mux_o_3737;
wire mux_o_3738;
wire mux_o_3739;
wire mux_o_3740;
wire mux_o_3741;
wire mux_o_3742;
wire mux_o_3743;
wire mux_o_3744;
wire mux_o_3745;
wire mux_o_3746;
wire mux_o_3747;
wire mux_o_3748;
wire mux_o_3749;
wire mux_o_3750;
wire mux_o_3751;
wire mux_o_3752;
wire mux_o_3753;
wire mux_o_3754;
wire mux_o_3755;
wire mux_o_3756;
wire mux_o_3757;
wire mux_o_3758;
wire mux_o_3759;
wire mux_o_3760;
wire mux_o_3761;
wire mux_o_3762;
wire mux_o_3763;
wire mux_o_3764;
wire mux_o_3765;
wire mux_o_3766;
wire mux_o_3767;
wire mux_o_3768;
wire mux_o_3769;
wire mux_o_3770;
wire mux_o_3771;
wire mux_o_3772;
wire mux_o_3773;
wire mux_o_3774;
wire mux_o_3775;
wire mux_o_3776;
wire mux_o_3777;
wire mux_o_3778;
wire mux_o_3779;
wire mux_o_3780;
wire mux_o_3781;
wire mux_o_3782;
wire mux_o_3783;
wire mux_o_3784;
wire mux_o_3785;
wire mux_o_3786;
wire mux_o_3787;
wire mux_o_3788;
wire mux_o_3789;
wire mux_o_3790;
wire mux_o_3791;
wire mux_o_3792;
wire mux_o_3793;
wire mux_o_3794;
wire mux_o_3795;
wire mux_o_3796;
wire mux_o_3797;
wire mux_o_3798;
wire mux_o_3799;
wire mux_o_3800;
wire mux_o_3801;
wire mux_o_3802;
wire mux_o_3803;
wire mux_o_3804;
wire mux_o_3805;
wire mux_o_3806;
wire mux_o_3807;
wire mux_o_3808;
wire mux_o_3810;
wire mux_o_3811;
wire mux_o_3812;
wire mux_o_3813;
wire mux_o_3814;
wire mux_o_3815;
wire mux_o_3816;
wire mux_o_3817;
wire mux_o_3818;
wire mux_o_3819;
wire mux_o_3820;
wire mux_o_3821;
wire mux_o_3822;
wire mux_o_3823;
wire mux_o_3824;
wire mux_o_3825;
wire mux_o_3826;
wire mux_o_3827;
wire mux_o_3828;
wire mux_o_3829;
wire mux_o_3830;
wire mux_o_3831;
wire mux_o_3832;
wire mux_o_3833;
wire mux_o_3834;
wire mux_o_3835;
wire mux_o_3836;
wire mux_o_3837;
wire mux_o_3838;
wire mux_o_3839;
wire mux_o_3840;
wire mux_o_3841;
wire mux_o_3842;
wire mux_o_3843;
wire mux_o_3844;
wire mux_o_3845;
wire mux_o_3846;
wire mux_o_3847;
wire mux_o_3848;
wire mux_o_3849;
wire mux_o_3850;
wire mux_o_3851;
wire mux_o_3852;
wire mux_o_3853;
wire mux_o_3854;
wire mux_o_3855;
wire mux_o_3856;
wire mux_o_3857;
wire mux_o_3858;
wire mux_o_3859;
wire mux_o_3860;
wire mux_o_3861;
wire mux_o_3862;
wire mux_o_3863;
wire mux_o_3864;
wire mux_o_3865;
wire mux_o_3866;
wire mux_o_3867;
wire mux_o_3868;
wire mux_o_3869;
wire mux_o_3870;
wire mux_o_3871;
wire mux_o_3872;
wire mux_o_3873;
wire mux_o_3874;
wire mux_o_3875;
wire mux_o_3876;
wire mux_o_3877;
wire mux_o_3878;
wire mux_o_3879;
wire mux_o_3880;
wire mux_o_3881;
wire mux_o_3882;
wire mux_o_3883;
wire mux_o_3884;
wire mux_o_3885;
wire mux_o_3886;
wire mux_o_3887;
wire mux_o_3888;
wire mux_o_3889;
wire mux_o_3890;
wire mux_o_3891;
wire mux_o_3892;
wire mux_o_3893;
wire mux_o_3894;
wire mux_o_3895;
wire mux_o_3896;
wire mux_o_3897;
wire mux_o_3898;
wire mux_o_3899;
wire mux_o_3900;
wire mux_o_3901;
wire mux_o_3902;
wire mux_o_3903;
wire mux_o_3904;
wire mux_o_3905;
wire mux_o_3906;
wire mux_o_3907;
wire mux_o_3908;
wire mux_o_3909;
wire mux_o_3910;
wire mux_o_3911;
wire mux_o_3912;
wire mux_o_3913;
wire mux_o_3914;
wire mux_o_3915;
wire mux_o_3916;
wire mux_o_3917;
wire mux_o_3918;
wire mux_o_3919;
wire mux_o_3920;
wire mux_o_3921;
wire mux_o_3922;
wire mux_o_3923;
wire mux_o_3924;
wire mux_o_3925;
wire mux_o_3926;
wire mux_o_3927;
wire mux_o_3928;
wire mux_o_3929;
wire mux_o_3930;
wire mux_o_3931;
wire mux_o_3932;
wire mux_o_3933;
wire mux_o_3934;
wire mux_o_3935;
wire mux_o_3937;
wire mux_o_3938;
wire mux_o_3939;
wire mux_o_3940;
wire mux_o_3941;
wire mux_o_3942;
wire mux_o_3943;
wire mux_o_3944;
wire mux_o_3945;
wire mux_o_3946;
wire mux_o_3947;
wire mux_o_3948;
wire mux_o_3949;
wire mux_o_3950;
wire mux_o_3951;
wire mux_o_3952;
wire mux_o_3953;
wire mux_o_3954;
wire mux_o_3955;
wire mux_o_3956;
wire mux_o_3957;
wire mux_o_3958;
wire mux_o_3959;
wire mux_o_3960;
wire mux_o_3961;
wire mux_o_3962;
wire mux_o_3963;
wire mux_o_3964;
wire mux_o_3965;
wire mux_o_3966;
wire mux_o_3967;
wire mux_o_3968;
wire mux_o_3969;
wire mux_o_3970;
wire mux_o_3971;
wire mux_o_3972;
wire mux_o_3973;
wire mux_o_3974;
wire mux_o_3975;
wire mux_o_3976;
wire mux_o_3977;
wire mux_o_3978;
wire mux_o_3979;
wire mux_o_3980;
wire mux_o_3981;
wire mux_o_3982;
wire mux_o_3983;
wire mux_o_3984;
wire mux_o_3985;
wire mux_o_3986;
wire mux_o_3987;
wire mux_o_3988;
wire mux_o_3989;
wire mux_o_3990;
wire mux_o_3991;
wire mux_o_3992;
wire mux_o_3993;
wire mux_o_3994;
wire mux_o_3995;
wire mux_o_3996;
wire mux_o_3997;
wire mux_o_3998;
wire mux_o_3999;
wire mux_o_4000;
wire mux_o_4001;
wire mux_o_4002;
wire mux_o_4003;
wire mux_o_4004;
wire mux_o_4005;
wire mux_o_4006;
wire mux_o_4007;
wire mux_o_4008;
wire mux_o_4009;
wire mux_o_4010;
wire mux_o_4011;
wire mux_o_4012;
wire mux_o_4013;
wire mux_o_4014;
wire mux_o_4015;
wire mux_o_4016;
wire mux_o_4017;
wire mux_o_4018;
wire mux_o_4019;
wire mux_o_4020;
wire mux_o_4021;
wire mux_o_4022;
wire mux_o_4023;
wire mux_o_4024;
wire mux_o_4025;
wire mux_o_4026;
wire mux_o_4027;
wire mux_o_4028;
wire mux_o_4029;
wire mux_o_4030;
wire mux_o_4031;
wire mux_o_4032;
wire mux_o_4033;
wire mux_o_4034;
wire mux_o_4035;
wire mux_o_4036;
wire mux_o_4037;
wire mux_o_4038;
wire mux_o_4039;
wire mux_o_4040;
wire mux_o_4041;
wire mux_o_4042;
wire mux_o_4043;
wire mux_o_4044;
wire mux_o_4045;
wire mux_o_4046;
wire mux_o_4047;
wire mux_o_4048;
wire mux_o_4049;
wire mux_o_4050;
wire mux_o_4051;
wire mux_o_4052;
wire mux_o_4053;
wire mux_o_4054;
wire mux_o_4055;
wire mux_o_4056;
wire mux_o_4057;
wire mux_o_4058;
wire mux_o_4059;
wire mux_o_4060;
wire mux_o_4061;
wire mux_o_4062;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT7 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_0.INIT = 128'h00000000000000000000000000000001;
LUT7 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_1.INIT = 128'h00000000000000000000000000000002;
LUT7 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_2.INIT = 128'h00000000000000000000000000000004;
LUT7 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_3.INIT = 128'h00000000000000000000000000000008;
LUT7 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_4.INIT = 128'h00000000000000000000000000000010;
LUT7 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_5.INIT = 128'h00000000000000000000000000000020;
LUT7 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_6.INIT = 128'h00000000000000000000000000000040;
LUT7 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_7.INIT = 128'h00000000000000000000000000000080;
LUT7 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_8.INIT = 128'h00000000000000000000000000000100;
LUT7 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_9.INIT = 128'h00000000000000000000000000000200;
LUT7 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_10.INIT = 128'h00000000000000000000000000000400;
LUT7 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_11.INIT = 128'h00000000000000000000000000000800;
LUT7 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_12.INIT = 128'h00000000000000000000000000001000;
LUT7 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_13.INIT = 128'h00000000000000000000000000002000;
LUT7 lut_inst_14 (
  .F(lut_f_14),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_14.INIT = 128'h00000000000000000000000000004000;
LUT7 lut_inst_15 (
  .F(lut_f_15),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_15.INIT = 128'h00000000000000000000000000008000;
LUT7 lut_inst_16 (
  .F(lut_f_16),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_16.INIT = 128'h00000000000000000000000000010000;
LUT7 lut_inst_17 (
  .F(lut_f_17),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_17.INIT = 128'h00000000000000000000000000020000;
LUT7 lut_inst_18 (
  .F(lut_f_18),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_18.INIT = 128'h00000000000000000000000000040000;
LUT7 lut_inst_19 (
  .F(lut_f_19),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_19.INIT = 128'h00000000000000000000000000080000;
LUT7 lut_inst_20 (
  .F(lut_f_20),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_20.INIT = 128'h00000000000000000000000000100000;
LUT7 lut_inst_21 (
  .F(lut_f_21),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_21.INIT = 128'h00000000000000000000000000200000;
LUT7 lut_inst_22 (
  .F(lut_f_22),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_22.INIT = 128'h00000000000000000000000000400000;
LUT7 lut_inst_23 (
  .F(lut_f_23),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_23.INIT = 128'h00000000000000000000000000800000;
LUT7 lut_inst_24 (
  .F(lut_f_24),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_24.INIT = 128'h00000000000000000000000001000000;
LUT7 lut_inst_25 (
  .F(lut_f_25),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_25.INIT = 128'h00000000000000000000000002000000;
LUT7 lut_inst_26 (
  .F(lut_f_26),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_26.INIT = 128'h00000000000000000000000004000000;
LUT7 lut_inst_27 (
  .F(lut_f_27),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_27.INIT = 128'h00000000000000000000000008000000;
LUT7 lut_inst_28 (
  .F(lut_f_28),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_28.INIT = 128'h00000000000000000000000010000000;
LUT7 lut_inst_29 (
  .F(lut_f_29),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_29.INIT = 128'h00000000000000000000000020000000;
LUT7 lut_inst_30 (
  .F(lut_f_30),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_30.INIT = 128'h00000000000000000000000040000000;
LUT7 lut_inst_31 (
  .F(lut_f_31),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_31.INIT = 128'h00000000000000000000000080000000;
LUT7 lut_inst_32 (
  .F(lut_f_32),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_32.INIT = 128'h00000000000000000000000100000000;
LUT7 lut_inst_33 (
  .F(lut_f_33),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_33.INIT = 128'h00000000000000000000000200000000;
LUT7 lut_inst_34 (
  .F(lut_f_34),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_34.INIT = 128'h00000000000000000000000400000000;
LUT7 lut_inst_35 (
  .F(lut_f_35),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_35.INIT = 128'h00000000000000000000000800000000;
LUT7 lut_inst_36 (
  .F(lut_f_36),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_36.INIT = 128'h00000000000000000000001000000000;
LUT7 lut_inst_37 (
  .F(lut_f_37),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_37.INIT = 128'h00000000000000000000002000000000;
LUT7 lut_inst_38 (
  .F(lut_f_38),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_38.INIT = 128'h00000000000000000000004000000000;
LUT7 lut_inst_39 (
  .F(lut_f_39),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_39.INIT = 128'h00000000000000000000008000000000;
LUT7 lut_inst_40 (
  .F(lut_f_40),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_40.INIT = 128'h00000000000000000000010000000000;
LUT7 lut_inst_41 (
  .F(lut_f_41),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_41.INIT = 128'h00000000000000000000020000000000;
LUT7 lut_inst_42 (
  .F(lut_f_42),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_42.INIT = 128'h00000000000000000000040000000000;
LUT7 lut_inst_43 (
  .F(lut_f_43),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_43.INIT = 128'h00000000000000000000080000000000;
LUT7 lut_inst_44 (
  .F(lut_f_44),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_44.INIT = 128'h00000000000000000000100000000000;
LUT7 lut_inst_45 (
  .F(lut_f_45),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_45.INIT = 128'h00000000000000000000200000000000;
LUT7 lut_inst_46 (
  .F(lut_f_46),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_46.INIT = 128'h00000000000000000000400000000000;
LUT7 lut_inst_47 (
  .F(lut_f_47),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_47.INIT = 128'h00000000000000000000800000000000;
LUT7 lut_inst_48 (
  .F(lut_f_48),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_48.INIT = 128'h00000000000000000001000000000000;
LUT7 lut_inst_49 (
  .F(lut_f_49),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_49.INIT = 128'h00000000000000000002000000000000;
LUT7 lut_inst_50 (
  .F(lut_f_50),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_50.INIT = 128'h00000000000000000004000000000000;
LUT7 lut_inst_51 (
  .F(lut_f_51),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_51.INIT = 128'h00000000000000000008000000000000;
LUT7 lut_inst_52 (
  .F(lut_f_52),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_52.INIT = 128'h00000000000000000010000000000000;
LUT7 lut_inst_53 (
  .F(lut_f_53),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_53.INIT = 128'h00000000000000000020000000000000;
LUT7 lut_inst_54 (
  .F(lut_f_54),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_54.INIT = 128'h00000000000000000040000000000000;
LUT7 lut_inst_55 (
  .F(lut_f_55),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_55.INIT = 128'h00000000000000000080000000000000;
LUT7 lut_inst_56 (
  .F(lut_f_56),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_56.INIT = 128'h00000000000000000100000000000000;
LUT7 lut_inst_57 (
  .F(lut_f_57),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_57.INIT = 128'h00000000000000000200000000000000;
LUT7 lut_inst_58 (
  .F(lut_f_58),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_58.INIT = 128'h00000000000000000400000000000000;
LUT7 lut_inst_59 (
  .F(lut_f_59),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_59.INIT = 128'h00000000000000000800000000000000;
LUT7 lut_inst_60 (
  .F(lut_f_60),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_60.INIT = 128'h00000000000000001000000000000000;
LUT7 lut_inst_61 (
  .F(lut_f_61),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_61.INIT = 128'h00000000000000002000000000000000;
LUT7 lut_inst_62 (
  .F(lut_f_62),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_62.INIT = 128'h00000000000000004000000000000000;
LUT7 lut_inst_63 (
  .F(lut_f_63),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_63.INIT = 128'h00000000000000008000000000000000;
LUT7 lut_inst_64 (
  .F(lut_f_64),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_64.INIT = 128'h00000000000000010000000000000000;
LUT7 lut_inst_65 (
  .F(lut_f_65),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_65.INIT = 128'h00000000000000020000000000000000;
LUT7 lut_inst_66 (
  .F(lut_f_66),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_66.INIT = 128'h00000000000000040000000000000000;
LUT7 lut_inst_67 (
  .F(lut_f_67),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_67.INIT = 128'h00000000000000080000000000000000;
LUT7 lut_inst_68 (
  .F(lut_f_68),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_68.INIT = 128'h00000000000000100000000000000000;
LUT7 lut_inst_69 (
  .F(lut_f_69),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_69.INIT = 128'h00000000000000200000000000000000;
LUT7 lut_inst_70 (
  .F(lut_f_70),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_70.INIT = 128'h00000000000000400000000000000000;
LUT7 lut_inst_71 (
  .F(lut_f_71),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_71.INIT = 128'h00000000000000800000000000000000;
LUT7 lut_inst_72 (
  .F(lut_f_72),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_72.INIT = 128'h00000000000001000000000000000000;
LUT7 lut_inst_73 (
  .F(lut_f_73),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_73.INIT = 128'h00000000000002000000000000000000;
LUT7 lut_inst_74 (
  .F(lut_f_74),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_74.INIT = 128'h00000000000004000000000000000000;
LUT7 lut_inst_75 (
  .F(lut_f_75),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_75.INIT = 128'h00000000000008000000000000000000;
LUT7 lut_inst_76 (
  .F(lut_f_76),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_76.INIT = 128'h00000000000010000000000000000000;
LUT7 lut_inst_77 (
  .F(lut_f_77),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_77.INIT = 128'h00000000000020000000000000000000;
LUT7 lut_inst_78 (
  .F(lut_f_78),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_78.INIT = 128'h00000000000040000000000000000000;
LUT7 lut_inst_79 (
  .F(lut_f_79),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_79.INIT = 128'h00000000000080000000000000000000;
LUT7 lut_inst_80 (
  .F(lut_f_80),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_80.INIT = 128'h00000000000100000000000000000000;
LUT7 lut_inst_81 (
  .F(lut_f_81),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_81.INIT = 128'h00000000000200000000000000000000;
LUT7 lut_inst_82 (
  .F(lut_f_82),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_82.INIT = 128'h00000000000400000000000000000000;
LUT7 lut_inst_83 (
  .F(lut_f_83),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_83.INIT = 128'h00000000000800000000000000000000;
LUT7 lut_inst_84 (
  .F(lut_f_84),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_84.INIT = 128'h00000000001000000000000000000000;
LUT7 lut_inst_85 (
  .F(lut_f_85),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_85.INIT = 128'h00000000002000000000000000000000;
LUT7 lut_inst_86 (
  .F(lut_f_86),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_86.INIT = 128'h00000000004000000000000000000000;
LUT7 lut_inst_87 (
  .F(lut_f_87),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_87.INIT = 128'h00000000008000000000000000000000;
LUT7 lut_inst_88 (
  .F(lut_f_88),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_88.INIT = 128'h00000000010000000000000000000000;
LUT7 lut_inst_89 (
  .F(lut_f_89),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_89.INIT = 128'h00000000020000000000000000000000;
LUT7 lut_inst_90 (
  .F(lut_f_90),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_90.INIT = 128'h00000000040000000000000000000000;
LUT7 lut_inst_91 (
  .F(lut_f_91),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_91.INIT = 128'h00000000080000000000000000000000;
LUT7 lut_inst_92 (
  .F(lut_f_92),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_92.INIT = 128'h00000000100000000000000000000000;
LUT7 lut_inst_93 (
  .F(lut_f_93),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_93.INIT = 128'h00000000200000000000000000000000;
LUT7 lut_inst_94 (
  .F(lut_f_94),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_94.INIT = 128'h00000000400000000000000000000000;
LUT7 lut_inst_95 (
  .F(lut_f_95),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_95.INIT = 128'h00000000800000000000000000000000;
LUT7 lut_inst_96 (
  .F(lut_f_96),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_96.INIT = 128'h00000001000000000000000000000000;
LUT7 lut_inst_97 (
  .F(lut_f_97),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_97.INIT = 128'h00000002000000000000000000000000;
LUT7 lut_inst_98 (
  .F(lut_f_98),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_98.INIT = 128'h00000004000000000000000000000000;
LUT7 lut_inst_99 (
  .F(lut_f_99),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_99.INIT = 128'h00000008000000000000000000000000;
LUT7 lut_inst_100 (
  .F(lut_f_100),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_100.INIT = 128'h00000010000000000000000000000000;
LUT7 lut_inst_101 (
  .F(lut_f_101),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_101.INIT = 128'h00000020000000000000000000000000;
LUT7 lut_inst_102 (
  .F(lut_f_102),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_102.INIT = 128'h00000040000000000000000000000000;
LUT7 lut_inst_103 (
  .F(lut_f_103),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_103.INIT = 128'h00000080000000000000000000000000;
LUT7 lut_inst_104 (
  .F(lut_f_104),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_104.INIT = 128'h00000100000000000000000000000000;
LUT7 lut_inst_105 (
  .F(lut_f_105),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_105.INIT = 128'h00000200000000000000000000000000;
LUT7 lut_inst_106 (
  .F(lut_f_106),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_106.INIT = 128'h00000400000000000000000000000000;
LUT7 lut_inst_107 (
  .F(lut_f_107),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_107.INIT = 128'h00000800000000000000000000000000;
LUT7 lut_inst_108 (
  .F(lut_f_108),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_108.INIT = 128'h00001000000000000000000000000000;
LUT7 lut_inst_109 (
  .F(lut_f_109),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_109.INIT = 128'h00002000000000000000000000000000;
LUT7 lut_inst_110 (
  .F(lut_f_110),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_110.INIT = 128'h00004000000000000000000000000000;
LUT7 lut_inst_111 (
  .F(lut_f_111),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_111.INIT = 128'h00008000000000000000000000000000;
LUT7 lut_inst_112 (
  .F(lut_f_112),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_112.INIT = 128'h00010000000000000000000000000000;
LUT7 lut_inst_113 (
  .F(lut_f_113),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_113.INIT = 128'h00020000000000000000000000000000;
LUT7 lut_inst_114 (
  .F(lut_f_114),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_114.INIT = 128'h00040000000000000000000000000000;
LUT7 lut_inst_115 (
  .F(lut_f_115),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_115.INIT = 128'h00080000000000000000000000000000;
LUT7 lut_inst_116 (
  .F(lut_f_116),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_116.INIT = 128'h00100000000000000000000000000000;
LUT7 lut_inst_117 (
  .F(lut_f_117),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_117.INIT = 128'h00200000000000000000000000000000;
LUT7 lut_inst_118 (
  .F(lut_f_118),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_118.INIT = 128'h00400000000000000000000000000000;
LUT7 lut_inst_119 (
  .F(lut_f_119),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_119.INIT = 128'h00800000000000000000000000000000;
LUT7 lut_inst_120 (
  .F(lut_f_120),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_120.INIT = 128'h01000000000000000000000000000000;
LUT7 lut_inst_121 (
  .F(lut_f_121),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_121.INIT = 128'h02000000000000000000000000000000;
LUT7 lut_inst_122 (
  .F(lut_f_122),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_122.INIT = 128'h04000000000000000000000000000000;
LUT7 lut_inst_123 (
  .F(lut_f_123),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_123.INIT = 128'h08000000000000000000000000000000;
LUT7 lut_inst_124 (
  .F(lut_f_124),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_124.INIT = 128'h10000000000000000000000000000000;
LUT7 lut_inst_125 (
  .F(lut_f_125),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_125.INIT = 128'h20000000000000000000000000000000;
LUT7 lut_inst_126 (
  .F(lut_f_126),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_126.INIT = 128'h40000000000000000000000000000000;
LUT7 lut_inst_127 (
  .F(lut_f_127),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_127.INIT = 128'h80000000000000000000000000000000;
LUT7 lut_inst_128 (
  .F(lut_f_128),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_128.INIT = 128'h00000000000000000000000000000001;
LUT7 lut_inst_129 (
  .F(lut_f_129),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_129.INIT = 128'h00000000000000000000000000000002;
LUT7 lut_inst_130 (
  .F(lut_f_130),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_130.INIT = 128'h00000000000000000000000000000004;
LUT7 lut_inst_131 (
  .F(lut_f_131),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_131.INIT = 128'h00000000000000000000000000000008;
LUT7 lut_inst_132 (
  .F(lut_f_132),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_132.INIT = 128'h00000000000000000000000000000010;
LUT7 lut_inst_133 (
  .F(lut_f_133),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_133.INIT = 128'h00000000000000000000000000000020;
LUT7 lut_inst_134 (
  .F(lut_f_134),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_134.INIT = 128'h00000000000000000000000000000040;
LUT7 lut_inst_135 (
  .F(lut_f_135),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_135.INIT = 128'h00000000000000000000000000000080;
LUT7 lut_inst_136 (
  .F(lut_f_136),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_136.INIT = 128'h00000000000000000000000000000100;
LUT7 lut_inst_137 (
  .F(lut_f_137),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_137.INIT = 128'h00000000000000000000000000000200;
LUT7 lut_inst_138 (
  .F(lut_f_138),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_138.INIT = 128'h00000000000000000000000000000400;
LUT7 lut_inst_139 (
  .F(lut_f_139),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_139.INIT = 128'h00000000000000000000000000000800;
LUT7 lut_inst_140 (
  .F(lut_f_140),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_140.INIT = 128'h00000000000000000000000000001000;
LUT7 lut_inst_141 (
  .F(lut_f_141),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_141.INIT = 128'h00000000000000000000000000002000;
LUT7 lut_inst_142 (
  .F(lut_f_142),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_142.INIT = 128'h00000000000000000000000000004000;
LUT7 lut_inst_143 (
  .F(lut_f_143),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_143.INIT = 128'h00000000000000000000000000008000;
LUT7 lut_inst_144 (
  .F(lut_f_144),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_144.INIT = 128'h00000000000000000000000000010000;
LUT7 lut_inst_145 (
  .F(lut_f_145),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_145.INIT = 128'h00000000000000000000000000020000;
LUT7 lut_inst_146 (
  .F(lut_f_146),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_146.INIT = 128'h00000000000000000000000000040000;
LUT7 lut_inst_147 (
  .F(lut_f_147),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_147.INIT = 128'h00000000000000000000000000080000;
LUT7 lut_inst_148 (
  .F(lut_f_148),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_148.INIT = 128'h00000000000000000000000000100000;
LUT7 lut_inst_149 (
  .F(lut_f_149),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_149.INIT = 128'h00000000000000000000000000200000;
LUT7 lut_inst_150 (
  .F(lut_f_150),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_150.INIT = 128'h00000000000000000000000000400000;
LUT7 lut_inst_151 (
  .F(lut_f_151),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_151.INIT = 128'h00000000000000000000000000800000;
LUT7 lut_inst_152 (
  .F(lut_f_152),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_152.INIT = 128'h00000000000000000000000001000000;
LUT7 lut_inst_153 (
  .F(lut_f_153),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_153.INIT = 128'h00000000000000000000000002000000;
LUT7 lut_inst_154 (
  .F(lut_f_154),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_154.INIT = 128'h00000000000000000000000004000000;
LUT7 lut_inst_155 (
  .F(lut_f_155),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_155.INIT = 128'h00000000000000000000000008000000;
LUT7 lut_inst_156 (
  .F(lut_f_156),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_156.INIT = 128'h00000000000000000000000010000000;
LUT7 lut_inst_157 (
  .F(lut_f_157),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_157.INIT = 128'h00000000000000000000000020000000;
LUT7 lut_inst_158 (
  .F(lut_f_158),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_158.INIT = 128'h00000000000000000000000040000000;
LUT7 lut_inst_159 (
  .F(lut_f_159),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_159.INIT = 128'h00000000000000000000000080000000;
LUT7 lut_inst_160 (
  .F(lut_f_160),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_160.INIT = 128'h00000000000000000000000100000000;
LUT7 lut_inst_161 (
  .F(lut_f_161),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_161.INIT = 128'h00000000000000000000000200000000;
LUT7 lut_inst_162 (
  .F(lut_f_162),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_162.INIT = 128'h00000000000000000000000400000000;
LUT7 lut_inst_163 (
  .F(lut_f_163),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_163.INIT = 128'h00000000000000000000000800000000;
LUT7 lut_inst_164 (
  .F(lut_f_164),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_164.INIT = 128'h00000000000000000000001000000000;
LUT7 lut_inst_165 (
  .F(lut_f_165),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_165.INIT = 128'h00000000000000000000002000000000;
LUT7 lut_inst_166 (
  .F(lut_f_166),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_166.INIT = 128'h00000000000000000000004000000000;
LUT7 lut_inst_167 (
  .F(lut_f_167),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_167.INIT = 128'h00000000000000000000008000000000;
LUT7 lut_inst_168 (
  .F(lut_f_168),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_168.INIT = 128'h00000000000000000000010000000000;
LUT7 lut_inst_169 (
  .F(lut_f_169),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_169.INIT = 128'h00000000000000000000020000000000;
LUT7 lut_inst_170 (
  .F(lut_f_170),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_170.INIT = 128'h00000000000000000000040000000000;
LUT7 lut_inst_171 (
  .F(lut_f_171),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_171.INIT = 128'h00000000000000000000080000000000;
LUT7 lut_inst_172 (
  .F(lut_f_172),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_172.INIT = 128'h00000000000000000000100000000000;
LUT7 lut_inst_173 (
  .F(lut_f_173),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_173.INIT = 128'h00000000000000000000200000000000;
LUT7 lut_inst_174 (
  .F(lut_f_174),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_174.INIT = 128'h00000000000000000000400000000000;
LUT7 lut_inst_175 (
  .F(lut_f_175),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_175.INIT = 128'h00000000000000000000800000000000;
LUT7 lut_inst_176 (
  .F(lut_f_176),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_176.INIT = 128'h00000000000000000001000000000000;
LUT7 lut_inst_177 (
  .F(lut_f_177),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_177.INIT = 128'h00000000000000000002000000000000;
LUT7 lut_inst_178 (
  .F(lut_f_178),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_178.INIT = 128'h00000000000000000004000000000000;
LUT7 lut_inst_179 (
  .F(lut_f_179),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_179.INIT = 128'h00000000000000000008000000000000;
LUT7 lut_inst_180 (
  .F(lut_f_180),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_180.INIT = 128'h00000000000000000010000000000000;
LUT7 lut_inst_181 (
  .F(lut_f_181),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_181.INIT = 128'h00000000000000000020000000000000;
LUT7 lut_inst_182 (
  .F(lut_f_182),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_182.INIT = 128'h00000000000000000040000000000000;
LUT7 lut_inst_183 (
  .F(lut_f_183),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_183.INIT = 128'h00000000000000000080000000000000;
LUT7 lut_inst_184 (
  .F(lut_f_184),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_184.INIT = 128'h00000000000000000100000000000000;
LUT7 lut_inst_185 (
  .F(lut_f_185),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_185.INIT = 128'h00000000000000000200000000000000;
LUT7 lut_inst_186 (
  .F(lut_f_186),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_186.INIT = 128'h00000000000000000400000000000000;
LUT7 lut_inst_187 (
  .F(lut_f_187),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_187.INIT = 128'h00000000000000000800000000000000;
LUT7 lut_inst_188 (
  .F(lut_f_188),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_188.INIT = 128'h00000000000000001000000000000000;
LUT7 lut_inst_189 (
  .F(lut_f_189),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_189.INIT = 128'h00000000000000002000000000000000;
LUT7 lut_inst_190 (
  .F(lut_f_190),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_190.INIT = 128'h00000000000000004000000000000000;
LUT7 lut_inst_191 (
  .F(lut_f_191),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_191.INIT = 128'h00000000000000008000000000000000;
LUT7 lut_inst_192 (
  .F(lut_f_192),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_192.INIT = 128'h00000000000000010000000000000000;
LUT7 lut_inst_193 (
  .F(lut_f_193),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_193.INIT = 128'h00000000000000020000000000000000;
LUT7 lut_inst_194 (
  .F(lut_f_194),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_194.INIT = 128'h00000000000000040000000000000000;
LUT7 lut_inst_195 (
  .F(lut_f_195),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_195.INIT = 128'h00000000000000080000000000000000;
LUT7 lut_inst_196 (
  .F(lut_f_196),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_196.INIT = 128'h00000000000000100000000000000000;
LUT7 lut_inst_197 (
  .F(lut_f_197),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_197.INIT = 128'h00000000000000200000000000000000;
LUT7 lut_inst_198 (
  .F(lut_f_198),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_198.INIT = 128'h00000000000000400000000000000000;
LUT7 lut_inst_199 (
  .F(lut_f_199),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_199.INIT = 128'h00000000000000800000000000000000;
LUT7 lut_inst_200 (
  .F(lut_f_200),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_200.INIT = 128'h00000000000001000000000000000000;
LUT7 lut_inst_201 (
  .F(lut_f_201),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_201.INIT = 128'h00000000000002000000000000000000;
LUT7 lut_inst_202 (
  .F(lut_f_202),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_202.INIT = 128'h00000000000004000000000000000000;
LUT7 lut_inst_203 (
  .F(lut_f_203),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_203.INIT = 128'h00000000000008000000000000000000;
LUT7 lut_inst_204 (
  .F(lut_f_204),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_204.INIT = 128'h00000000000010000000000000000000;
LUT7 lut_inst_205 (
  .F(lut_f_205),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_205.INIT = 128'h00000000000020000000000000000000;
LUT7 lut_inst_206 (
  .F(lut_f_206),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_206.INIT = 128'h00000000000040000000000000000000;
LUT7 lut_inst_207 (
  .F(lut_f_207),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_207.INIT = 128'h00000000000080000000000000000000;
LUT7 lut_inst_208 (
  .F(lut_f_208),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_208.INIT = 128'h00000000000100000000000000000000;
LUT7 lut_inst_209 (
  .F(lut_f_209),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_209.INIT = 128'h00000000000200000000000000000000;
LUT7 lut_inst_210 (
  .F(lut_f_210),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_210.INIT = 128'h00000000000400000000000000000000;
LUT7 lut_inst_211 (
  .F(lut_f_211),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_211.INIT = 128'h00000000000800000000000000000000;
LUT7 lut_inst_212 (
  .F(lut_f_212),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_212.INIT = 128'h00000000001000000000000000000000;
LUT7 lut_inst_213 (
  .F(lut_f_213),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_213.INIT = 128'h00000000002000000000000000000000;
LUT7 lut_inst_214 (
  .F(lut_f_214),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_214.INIT = 128'h00000000004000000000000000000000;
LUT7 lut_inst_215 (
  .F(lut_f_215),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_215.INIT = 128'h00000000008000000000000000000000;
LUT7 lut_inst_216 (
  .F(lut_f_216),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_216.INIT = 128'h00000000010000000000000000000000;
LUT7 lut_inst_217 (
  .F(lut_f_217),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_217.INIT = 128'h00000000020000000000000000000000;
LUT7 lut_inst_218 (
  .F(lut_f_218),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_218.INIT = 128'h00000000040000000000000000000000;
LUT7 lut_inst_219 (
  .F(lut_f_219),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_219.INIT = 128'h00000000080000000000000000000000;
LUT7 lut_inst_220 (
  .F(lut_f_220),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_220.INIT = 128'h00000000100000000000000000000000;
LUT7 lut_inst_221 (
  .F(lut_f_221),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_221.INIT = 128'h00000000200000000000000000000000;
LUT7 lut_inst_222 (
  .F(lut_f_222),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_222.INIT = 128'h00000000400000000000000000000000;
LUT7 lut_inst_223 (
  .F(lut_f_223),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_223.INIT = 128'h00000000800000000000000000000000;
LUT7 lut_inst_224 (
  .F(lut_f_224),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_224.INIT = 128'h00000001000000000000000000000000;
LUT7 lut_inst_225 (
  .F(lut_f_225),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_225.INIT = 128'h00000002000000000000000000000000;
LUT7 lut_inst_226 (
  .F(lut_f_226),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_226.INIT = 128'h00000004000000000000000000000000;
LUT7 lut_inst_227 (
  .F(lut_f_227),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_227.INIT = 128'h00000008000000000000000000000000;
LUT7 lut_inst_228 (
  .F(lut_f_228),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_228.INIT = 128'h00000010000000000000000000000000;
LUT7 lut_inst_229 (
  .F(lut_f_229),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_229.INIT = 128'h00000020000000000000000000000000;
LUT7 lut_inst_230 (
  .F(lut_f_230),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_230.INIT = 128'h00000040000000000000000000000000;
LUT7 lut_inst_231 (
  .F(lut_f_231),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_231.INIT = 128'h00000080000000000000000000000000;
LUT7 lut_inst_232 (
  .F(lut_f_232),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_232.INIT = 128'h00000100000000000000000000000000;
LUT7 lut_inst_233 (
  .F(lut_f_233),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_233.INIT = 128'h00000200000000000000000000000000;
LUT7 lut_inst_234 (
  .F(lut_f_234),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_234.INIT = 128'h00000400000000000000000000000000;
LUT7 lut_inst_235 (
  .F(lut_f_235),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_235.INIT = 128'h00000800000000000000000000000000;
LUT7 lut_inst_236 (
  .F(lut_f_236),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_236.INIT = 128'h00001000000000000000000000000000;
LUT7 lut_inst_237 (
  .F(lut_f_237),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_237.INIT = 128'h00002000000000000000000000000000;
LUT7 lut_inst_238 (
  .F(lut_f_238),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_238.INIT = 128'h00004000000000000000000000000000;
LUT7 lut_inst_239 (
  .F(lut_f_239),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_239.INIT = 128'h00008000000000000000000000000000;
LUT7 lut_inst_240 (
  .F(lut_f_240),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_240.INIT = 128'h00010000000000000000000000000000;
LUT7 lut_inst_241 (
  .F(lut_f_241),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_241.INIT = 128'h00020000000000000000000000000000;
LUT7 lut_inst_242 (
  .F(lut_f_242),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_242.INIT = 128'h00040000000000000000000000000000;
LUT7 lut_inst_243 (
  .F(lut_f_243),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_243.INIT = 128'h00080000000000000000000000000000;
LUT7 lut_inst_244 (
  .F(lut_f_244),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_244.INIT = 128'h00100000000000000000000000000000;
LUT7 lut_inst_245 (
  .F(lut_f_245),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_245.INIT = 128'h00200000000000000000000000000000;
LUT7 lut_inst_246 (
  .F(lut_f_246),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_246.INIT = 128'h00400000000000000000000000000000;
LUT7 lut_inst_247 (
  .F(lut_f_247),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_247.INIT = 128'h00800000000000000000000000000000;
LUT7 lut_inst_248 (
  .F(lut_f_248),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_248.INIT = 128'h01000000000000000000000000000000;
LUT7 lut_inst_249 (
  .F(lut_f_249),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_249.INIT = 128'h02000000000000000000000000000000;
LUT7 lut_inst_250 (
  .F(lut_f_250),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_250.INIT = 128'h04000000000000000000000000000000;
LUT7 lut_inst_251 (
  .F(lut_f_251),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_251.INIT = 128'h08000000000000000000000000000000;
LUT7 lut_inst_252 (
  .F(lut_f_252),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_252.INIT = 128'h10000000000000000000000000000000;
LUT7 lut_inst_253 (
  .F(lut_f_253),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_253.INIT = 128'h20000000000000000000000000000000;
LUT7 lut_inst_254 (
  .F(lut_f_254),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_254.INIT = 128'h40000000000000000000000000000000;
LUT7 lut_inst_255 (
  .F(lut_f_255),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_255.INIT = 128'h80000000000000000000000000000000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],sdpb_inst_0_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_128}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_0.RESET_MODE = "SYNC";

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[15:0],sdpb_inst_1_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_129}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 16;
defparam sdpb_inst_1.BIT_WIDTH_1 = 16;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[15:0],sdpb_inst_2_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_130}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 16;
defparam sdpb_inst_2.BIT_WIDTH_1 = 16;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_2.RESET_MODE = "SYNC";

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[15:0],sdpb_inst_3_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_131}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 16;
defparam sdpb_inst_3.BIT_WIDTH_1 = 16;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[15:0],sdpb_inst_4_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_132}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 16;
defparam sdpb_inst_4.BIT_WIDTH_1 = 16;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_4.RESET_MODE = "SYNC";

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[15:0],sdpb_inst_5_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_133}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 16;
defparam sdpb_inst_5.BIT_WIDTH_1 = 16;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[15:0],sdpb_inst_6_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_134}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 16;
defparam sdpb_inst_6.BIT_WIDTH_1 = 16;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_6.RESET_MODE = "SYNC";

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[15:0],sdpb_inst_7_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_135}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 16;
defparam sdpb_inst_7.BIT_WIDTH_1 = 16;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[15:0],sdpb_inst_8_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_136}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 16;
defparam sdpb_inst_8.BIT_WIDTH_1 = 16;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[15:0],sdpb_inst_9_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_137}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_9.READ_MODE = 1'b0;
defparam sdpb_inst_9.BIT_WIDTH_0 = 16;
defparam sdpb_inst_9.BIT_WIDTH_1 = 16;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_9.RESET_MODE = "SYNC";

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[15:0],sdpb_inst_10_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_138}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_10.READ_MODE = 1'b0;
defparam sdpb_inst_10.BIT_WIDTH_0 = 16;
defparam sdpb_inst_10.BIT_WIDTH_1 = 16;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_10.RESET_MODE = "SYNC";

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[15:0],sdpb_inst_11_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_139}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_11.READ_MODE = 1'b0;
defparam sdpb_inst_11.BIT_WIDTH_0 = 16;
defparam sdpb_inst_11.BIT_WIDTH_1 = 16;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_11.RESET_MODE = "SYNC";

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[15:0],sdpb_inst_12_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_140}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_12.READ_MODE = 1'b0;
defparam sdpb_inst_12.BIT_WIDTH_0 = 16;
defparam sdpb_inst_12.BIT_WIDTH_1 = 16;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_12.RESET_MODE = "SYNC";

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[15:0],sdpb_inst_13_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_141}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_13.READ_MODE = 1'b0;
defparam sdpb_inst_13.BIT_WIDTH_0 = 16;
defparam sdpb_inst_13.BIT_WIDTH_1 = 16;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_13.RESET_MODE = "SYNC";

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[15:0],sdpb_inst_14_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_142}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_14.READ_MODE = 1'b0;
defparam sdpb_inst_14.BIT_WIDTH_0 = 16;
defparam sdpb_inst_14.BIT_WIDTH_1 = 16;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_14.RESET_MODE = "SYNC";

SDPB sdpb_inst_15 (
    .DO({sdpb_inst_15_dout_w[15:0],sdpb_inst_15_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_143}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_15.READ_MODE = 1'b0;
defparam sdpb_inst_15.BIT_WIDTH_0 = 16;
defparam sdpb_inst_15.BIT_WIDTH_1 = 16;
defparam sdpb_inst_15.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_15.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_15.RESET_MODE = "SYNC";

SDPB sdpb_inst_16 (
    .DO({sdpb_inst_16_dout_w[15:0],sdpb_inst_16_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_16}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_144}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_16.READ_MODE = 1'b0;
defparam sdpb_inst_16.BIT_WIDTH_0 = 16;
defparam sdpb_inst_16.BIT_WIDTH_1 = 16;
defparam sdpb_inst_16.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_16.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_16.RESET_MODE = "SYNC";

SDPB sdpb_inst_17 (
    .DO({sdpb_inst_17_dout_w[15:0],sdpb_inst_17_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_17}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_145}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_17.READ_MODE = 1'b0;
defparam sdpb_inst_17.BIT_WIDTH_0 = 16;
defparam sdpb_inst_17.BIT_WIDTH_1 = 16;
defparam sdpb_inst_17.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_17.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_17.RESET_MODE = "SYNC";

SDPB sdpb_inst_18 (
    .DO({sdpb_inst_18_dout_w[15:0],sdpb_inst_18_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_18}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_146}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_18.READ_MODE = 1'b0;
defparam sdpb_inst_18.BIT_WIDTH_0 = 16;
defparam sdpb_inst_18.BIT_WIDTH_1 = 16;
defparam sdpb_inst_18.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_18.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_18.RESET_MODE = "SYNC";

SDPB sdpb_inst_19 (
    .DO({sdpb_inst_19_dout_w[15:0],sdpb_inst_19_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_19}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_147}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_19.READ_MODE = 1'b0;
defparam sdpb_inst_19.BIT_WIDTH_0 = 16;
defparam sdpb_inst_19.BIT_WIDTH_1 = 16;
defparam sdpb_inst_19.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_19.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_19.RESET_MODE = "SYNC";

SDPB sdpb_inst_20 (
    .DO({sdpb_inst_20_dout_w[15:0],sdpb_inst_20_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_20}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_148}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_20.READ_MODE = 1'b0;
defparam sdpb_inst_20.BIT_WIDTH_0 = 16;
defparam sdpb_inst_20.BIT_WIDTH_1 = 16;
defparam sdpb_inst_20.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_20.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_20.RESET_MODE = "SYNC";

SDPB sdpb_inst_21 (
    .DO({sdpb_inst_21_dout_w[15:0],sdpb_inst_21_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_21}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_149}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_21.READ_MODE = 1'b0;
defparam sdpb_inst_21.BIT_WIDTH_0 = 16;
defparam sdpb_inst_21.BIT_WIDTH_1 = 16;
defparam sdpb_inst_21.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_21.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_21.RESET_MODE = "SYNC";

SDPB sdpb_inst_22 (
    .DO({sdpb_inst_22_dout_w[15:0],sdpb_inst_22_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_22}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_150}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_22.READ_MODE = 1'b0;
defparam sdpb_inst_22.BIT_WIDTH_0 = 16;
defparam sdpb_inst_22.BIT_WIDTH_1 = 16;
defparam sdpb_inst_22.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_22.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_22.RESET_MODE = "SYNC";

SDPB sdpb_inst_23 (
    .DO({sdpb_inst_23_dout_w[15:0],sdpb_inst_23_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_23}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_151}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_23.READ_MODE = 1'b0;
defparam sdpb_inst_23.BIT_WIDTH_0 = 16;
defparam sdpb_inst_23.BIT_WIDTH_1 = 16;
defparam sdpb_inst_23.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_23.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_23.RESET_MODE = "SYNC";

SDPB sdpb_inst_24 (
    .DO({sdpb_inst_24_dout_w[15:0],sdpb_inst_24_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_24}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_152}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_24.READ_MODE = 1'b0;
defparam sdpb_inst_24.BIT_WIDTH_0 = 16;
defparam sdpb_inst_24.BIT_WIDTH_1 = 16;
defparam sdpb_inst_24.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_24.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_24.RESET_MODE = "SYNC";

SDPB sdpb_inst_25 (
    .DO({sdpb_inst_25_dout_w[15:0],sdpb_inst_25_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_25}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_153}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_25.READ_MODE = 1'b0;
defparam sdpb_inst_25.BIT_WIDTH_0 = 16;
defparam sdpb_inst_25.BIT_WIDTH_1 = 16;
defparam sdpb_inst_25.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_25.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_25.RESET_MODE = "SYNC";

SDPB sdpb_inst_26 (
    .DO({sdpb_inst_26_dout_w[15:0],sdpb_inst_26_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_26}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_154}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_26.READ_MODE = 1'b0;
defparam sdpb_inst_26.BIT_WIDTH_0 = 16;
defparam sdpb_inst_26.BIT_WIDTH_1 = 16;
defparam sdpb_inst_26.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_26.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_26.RESET_MODE = "SYNC";

SDPB sdpb_inst_27 (
    .DO({sdpb_inst_27_dout_w[15:0],sdpb_inst_27_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_27}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_155}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_27.READ_MODE = 1'b0;
defparam sdpb_inst_27.BIT_WIDTH_0 = 16;
defparam sdpb_inst_27.BIT_WIDTH_1 = 16;
defparam sdpb_inst_27.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_27.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_27.RESET_MODE = "SYNC";

SDPB sdpb_inst_28 (
    .DO({sdpb_inst_28_dout_w[15:0],sdpb_inst_28_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_28}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_156}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_28.READ_MODE = 1'b0;
defparam sdpb_inst_28.BIT_WIDTH_0 = 16;
defparam sdpb_inst_28.BIT_WIDTH_1 = 16;
defparam sdpb_inst_28.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_28.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_28.RESET_MODE = "SYNC";

SDPB sdpb_inst_29 (
    .DO({sdpb_inst_29_dout_w[15:0],sdpb_inst_29_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_29}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_157}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_29.READ_MODE = 1'b0;
defparam sdpb_inst_29.BIT_WIDTH_0 = 16;
defparam sdpb_inst_29.BIT_WIDTH_1 = 16;
defparam sdpb_inst_29.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_29.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_29.RESET_MODE = "SYNC";

SDPB sdpb_inst_30 (
    .DO({sdpb_inst_30_dout_w[15:0],sdpb_inst_30_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_30}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_158}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_30.READ_MODE = 1'b0;
defparam sdpb_inst_30.BIT_WIDTH_0 = 16;
defparam sdpb_inst_30.BIT_WIDTH_1 = 16;
defparam sdpb_inst_30.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_30.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_30.RESET_MODE = "SYNC";

SDPB sdpb_inst_31 (
    .DO({sdpb_inst_31_dout_w[15:0],sdpb_inst_31_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_31}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_159}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_31.READ_MODE = 1'b0;
defparam sdpb_inst_31.BIT_WIDTH_0 = 16;
defparam sdpb_inst_31.BIT_WIDTH_1 = 16;
defparam sdpb_inst_31.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_31.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_31.RESET_MODE = "SYNC";

SDPB sdpb_inst_32 (
    .DO({sdpb_inst_32_dout_w[15:0],sdpb_inst_32_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_32}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_160}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_32.READ_MODE = 1'b0;
defparam sdpb_inst_32.BIT_WIDTH_0 = 16;
defparam sdpb_inst_32.BIT_WIDTH_1 = 16;
defparam sdpb_inst_32.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_32.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_32.RESET_MODE = "SYNC";

SDPB sdpb_inst_33 (
    .DO({sdpb_inst_33_dout_w[15:0],sdpb_inst_33_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_33}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_161}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_33.READ_MODE = 1'b0;
defparam sdpb_inst_33.BIT_WIDTH_0 = 16;
defparam sdpb_inst_33.BIT_WIDTH_1 = 16;
defparam sdpb_inst_33.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_33.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_33.RESET_MODE = "SYNC";

SDPB sdpb_inst_34 (
    .DO({sdpb_inst_34_dout_w[15:0],sdpb_inst_34_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_34}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_162}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_34.READ_MODE = 1'b0;
defparam sdpb_inst_34.BIT_WIDTH_0 = 16;
defparam sdpb_inst_34.BIT_WIDTH_1 = 16;
defparam sdpb_inst_34.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_34.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_34.RESET_MODE = "SYNC";

SDPB sdpb_inst_35 (
    .DO({sdpb_inst_35_dout_w[15:0],sdpb_inst_35_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_35}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_163}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_35.READ_MODE = 1'b0;
defparam sdpb_inst_35.BIT_WIDTH_0 = 16;
defparam sdpb_inst_35.BIT_WIDTH_1 = 16;
defparam sdpb_inst_35.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_35.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_35.RESET_MODE = "SYNC";

SDPB sdpb_inst_36 (
    .DO({sdpb_inst_36_dout_w[15:0],sdpb_inst_36_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_36}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_164}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_36.READ_MODE = 1'b0;
defparam sdpb_inst_36.BIT_WIDTH_0 = 16;
defparam sdpb_inst_36.BIT_WIDTH_1 = 16;
defparam sdpb_inst_36.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_36.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_36.RESET_MODE = "SYNC";

SDPB sdpb_inst_37 (
    .DO({sdpb_inst_37_dout_w[15:0],sdpb_inst_37_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_37}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_165}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_37.READ_MODE = 1'b0;
defparam sdpb_inst_37.BIT_WIDTH_0 = 16;
defparam sdpb_inst_37.BIT_WIDTH_1 = 16;
defparam sdpb_inst_37.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_37.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_37.RESET_MODE = "SYNC";

SDPB sdpb_inst_38 (
    .DO({sdpb_inst_38_dout_w[15:0],sdpb_inst_38_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_38}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_166}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_38.READ_MODE = 1'b0;
defparam sdpb_inst_38.BIT_WIDTH_0 = 16;
defparam sdpb_inst_38.BIT_WIDTH_1 = 16;
defparam sdpb_inst_38.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_38.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_38.RESET_MODE = "SYNC";

SDPB sdpb_inst_39 (
    .DO({sdpb_inst_39_dout_w[15:0],sdpb_inst_39_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_39}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_167}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_39.READ_MODE = 1'b0;
defparam sdpb_inst_39.BIT_WIDTH_0 = 16;
defparam sdpb_inst_39.BIT_WIDTH_1 = 16;
defparam sdpb_inst_39.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_39.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_39.RESET_MODE = "SYNC";

SDPB sdpb_inst_40 (
    .DO({sdpb_inst_40_dout_w[15:0],sdpb_inst_40_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_40}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_168}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_40.READ_MODE = 1'b0;
defparam sdpb_inst_40.BIT_WIDTH_0 = 16;
defparam sdpb_inst_40.BIT_WIDTH_1 = 16;
defparam sdpb_inst_40.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_40.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_40.RESET_MODE = "SYNC";

SDPB sdpb_inst_41 (
    .DO({sdpb_inst_41_dout_w[15:0],sdpb_inst_41_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_41}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_169}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_41.READ_MODE = 1'b0;
defparam sdpb_inst_41.BIT_WIDTH_0 = 16;
defparam sdpb_inst_41.BIT_WIDTH_1 = 16;
defparam sdpb_inst_41.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_41.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_41.RESET_MODE = "SYNC";

SDPB sdpb_inst_42 (
    .DO({sdpb_inst_42_dout_w[15:0],sdpb_inst_42_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_42}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_170}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_42.READ_MODE = 1'b0;
defparam sdpb_inst_42.BIT_WIDTH_0 = 16;
defparam sdpb_inst_42.BIT_WIDTH_1 = 16;
defparam sdpb_inst_42.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_42.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_42.RESET_MODE = "SYNC";

SDPB sdpb_inst_43 (
    .DO({sdpb_inst_43_dout_w[15:0],sdpb_inst_43_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_43}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_171}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_43.READ_MODE = 1'b0;
defparam sdpb_inst_43.BIT_WIDTH_0 = 16;
defparam sdpb_inst_43.BIT_WIDTH_1 = 16;
defparam sdpb_inst_43.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_43.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_43.RESET_MODE = "SYNC";

SDPB sdpb_inst_44 (
    .DO({sdpb_inst_44_dout_w[15:0],sdpb_inst_44_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_44}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_172}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_44.READ_MODE = 1'b0;
defparam sdpb_inst_44.BIT_WIDTH_0 = 16;
defparam sdpb_inst_44.BIT_WIDTH_1 = 16;
defparam sdpb_inst_44.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_44.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_44.RESET_MODE = "SYNC";

SDPB sdpb_inst_45 (
    .DO({sdpb_inst_45_dout_w[15:0],sdpb_inst_45_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_45}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_173}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_45.READ_MODE = 1'b0;
defparam sdpb_inst_45.BIT_WIDTH_0 = 16;
defparam sdpb_inst_45.BIT_WIDTH_1 = 16;
defparam sdpb_inst_45.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_45.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_45.RESET_MODE = "SYNC";

SDPB sdpb_inst_46 (
    .DO({sdpb_inst_46_dout_w[15:0],sdpb_inst_46_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_46}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_174}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_46.READ_MODE = 1'b0;
defparam sdpb_inst_46.BIT_WIDTH_0 = 16;
defparam sdpb_inst_46.BIT_WIDTH_1 = 16;
defparam sdpb_inst_46.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_46.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_46.RESET_MODE = "SYNC";

SDPB sdpb_inst_47 (
    .DO({sdpb_inst_47_dout_w[15:0],sdpb_inst_47_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_47}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_175}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_47.READ_MODE = 1'b0;
defparam sdpb_inst_47.BIT_WIDTH_0 = 16;
defparam sdpb_inst_47.BIT_WIDTH_1 = 16;
defparam sdpb_inst_47.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_47.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_47.RESET_MODE = "SYNC";

SDPB sdpb_inst_48 (
    .DO({sdpb_inst_48_dout_w[15:0],sdpb_inst_48_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_48}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_176}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_48.READ_MODE = 1'b0;
defparam sdpb_inst_48.BIT_WIDTH_0 = 16;
defparam sdpb_inst_48.BIT_WIDTH_1 = 16;
defparam sdpb_inst_48.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_48.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_48.RESET_MODE = "SYNC";

SDPB sdpb_inst_49 (
    .DO({sdpb_inst_49_dout_w[15:0],sdpb_inst_49_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_49}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_177}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_49.READ_MODE = 1'b0;
defparam sdpb_inst_49.BIT_WIDTH_0 = 16;
defparam sdpb_inst_49.BIT_WIDTH_1 = 16;
defparam sdpb_inst_49.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_49.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_49.RESET_MODE = "SYNC";

SDPB sdpb_inst_50 (
    .DO({sdpb_inst_50_dout_w[15:0],sdpb_inst_50_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_50}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_178}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_50.READ_MODE = 1'b0;
defparam sdpb_inst_50.BIT_WIDTH_0 = 16;
defparam sdpb_inst_50.BIT_WIDTH_1 = 16;
defparam sdpb_inst_50.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_50.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_50.RESET_MODE = "SYNC";

SDPB sdpb_inst_51 (
    .DO({sdpb_inst_51_dout_w[15:0],sdpb_inst_51_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_51}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_179}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_51.READ_MODE = 1'b0;
defparam sdpb_inst_51.BIT_WIDTH_0 = 16;
defparam sdpb_inst_51.BIT_WIDTH_1 = 16;
defparam sdpb_inst_51.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_51.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_51.RESET_MODE = "SYNC";

SDPB sdpb_inst_52 (
    .DO({sdpb_inst_52_dout_w[15:0],sdpb_inst_52_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_52}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_180}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_52.READ_MODE = 1'b0;
defparam sdpb_inst_52.BIT_WIDTH_0 = 16;
defparam sdpb_inst_52.BIT_WIDTH_1 = 16;
defparam sdpb_inst_52.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_52.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_52.RESET_MODE = "SYNC";

SDPB sdpb_inst_53 (
    .DO({sdpb_inst_53_dout_w[15:0],sdpb_inst_53_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_53}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_181}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_53.READ_MODE = 1'b0;
defparam sdpb_inst_53.BIT_WIDTH_0 = 16;
defparam sdpb_inst_53.BIT_WIDTH_1 = 16;
defparam sdpb_inst_53.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_53.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_53.RESET_MODE = "SYNC";

SDPB sdpb_inst_54 (
    .DO({sdpb_inst_54_dout_w[15:0],sdpb_inst_54_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_54}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_182}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_54.READ_MODE = 1'b0;
defparam sdpb_inst_54.BIT_WIDTH_0 = 16;
defparam sdpb_inst_54.BIT_WIDTH_1 = 16;
defparam sdpb_inst_54.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_54.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_54.RESET_MODE = "SYNC";

SDPB sdpb_inst_55 (
    .DO({sdpb_inst_55_dout_w[15:0],sdpb_inst_55_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_55}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_183}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_55.READ_MODE = 1'b0;
defparam sdpb_inst_55.BIT_WIDTH_0 = 16;
defparam sdpb_inst_55.BIT_WIDTH_1 = 16;
defparam sdpb_inst_55.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_55.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_55.RESET_MODE = "SYNC";

SDPB sdpb_inst_56 (
    .DO({sdpb_inst_56_dout_w[15:0],sdpb_inst_56_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_184}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_56.READ_MODE = 1'b0;
defparam sdpb_inst_56.BIT_WIDTH_0 = 16;
defparam sdpb_inst_56.BIT_WIDTH_1 = 16;
defparam sdpb_inst_56.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_56.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_56.RESET_MODE = "SYNC";

SDPB sdpb_inst_57 (
    .DO({sdpb_inst_57_dout_w[15:0],sdpb_inst_57_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_185}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_57.READ_MODE = 1'b0;
defparam sdpb_inst_57.BIT_WIDTH_0 = 16;
defparam sdpb_inst_57.BIT_WIDTH_1 = 16;
defparam sdpb_inst_57.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_57.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_57.RESET_MODE = "SYNC";

SDPB sdpb_inst_58 (
    .DO({sdpb_inst_58_dout_w[15:0],sdpb_inst_58_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_58}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_186}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_58.READ_MODE = 1'b0;
defparam sdpb_inst_58.BIT_WIDTH_0 = 16;
defparam sdpb_inst_58.BIT_WIDTH_1 = 16;
defparam sdpb_inst_58.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_58.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_58.RESET_MODE = "SYNC";

SDPB sdpb_inst_59 (
    .DO({sdpb_inst_59_dout_w[15:0],sdpb_inst_59_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_59}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_187}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_59.READ_MODE = 1'b0;
defparam sdpb_inst_59.BIT_WIDTH_0 = 16;
defparam sdpb_inst_59.BIT_WIDTH_1 = 16;
defparam sdpb_inst_59.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_59.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_59.RESET_MODE = "SYNC";

SDPB sdpb_inst_60 (
    .DO({sdpb_inst_60_dout_w[15:0],sdpb_inst_60_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_60}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_188}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_60.READ_MODE = 1'b0;
defparam sdpb_inst_60.BIT_WIDTH_0 = 16;
defparam sdpb_inst_60.BIT_WIDTH_1 = 16;
defparam sdpb_inst_60.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_60.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_60.RESET_MODE = "SYNC";

SDPB sdpb_inst_61 (
    .DO({sdpb_inst_61_dout_w[15:0],sdpb_inst_61_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_61}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_189}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_61.READ_MODE = 1'b0;
defparam sdpb_inst_61.BIT_WIDTH_0 = 16;
defparam sdpb_inst_61.BIT_WIDTH_1 = 16;
defparam sdpb_inst_61.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_61.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_61.RESET_MODE = "SYNC";

SDPB sdpb_inst_62 (
    .DO({sdpb_inst_62_dout_w[15:0],sdpb_inst_62_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_62}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_190}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_62.READ_MODE = 1'b0;
defparam sdpb_inst_62.BIT_WIDTH_0 = 16;
defparam sdpb_inst_62.BIT_WIDTH_1 = 16;
defparam sdpb_inst_62.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_62.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_62.RESET_MODE = "SYNC";

SDPB sdpb_inst_63 (
    .DO({sdpb_inst_63_dout_w[15:0],sdpb_inst_63_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_63}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_191}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_63.READ_MODE = 1'b0;
defparam sdpb_inst_63.BIT_WIDTH_0 = 16;
defparam sdpb_inst_63.BIT_WIDTH_1 = 16;
defparam sdpb_inst_63.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_63.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_63.RESET_MODE = "SYNC";

SDPB sdpb_inst_64 (
    .DO({sdpb_inst_64_dout_w[15:0],sdpb_inst_64_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_64}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_192}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_64.READ_MODE = 1'b0;
defparam sdpb_inst_64.BIT_WIDTH_0 = 16;
defparam sdpb_inst_64.BIT_WIDTH_1 = 16;
defparam sdpb_inst_64.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_64.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_64.RESET_MODE = "SYNC";

SDPB sdpb_inst_65 (
    .DO({sdpb_inst_65_dout_w[15:0],sdpb_inst_65_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_65}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_193}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_65.READ_MODE = 1'b0;
defparam sdpb_inst_65.BIT_WIDTH_0 = 16;
defparam sdpb_inst_65.BIT_WIDTH_1 = 16;
defparam sdpb_inst_65.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_65.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_65.RESET_MODE = "SYNC";

SDPB sdpb_inst_66 (
    .DO({sdpb_inst_66_dout_w[15:0],sdpb_inst_66_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_66}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_194}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_66.READ_MODE = 1'b0;
defparam sdpb_inst_66.BIT_WIDTH_0 = 16;
defparam sdpb_inst_66.BIT_WIDTH_1 = 16;
defparam sdpb_inst_66.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_66.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_66.RESET_MODE = "SYNC";

SDPB sdpb_inst_67 (
    .DO({sdpb_inst_67_dout_w[15:0],sdpb_inst_67_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_67}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_195}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_67.READ_MODE = 1'b0;
defparam sdpb_inst_67.BIT_WIDTH_0 = 16;
defparam sdpb_inst_67.BIT_WIDTH_1 = 16;
defparam sdpb_inst_67.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_67.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_67.RESET_MODE = "SYNC";

SDPB sdpb_inst_68 (
    .DO({sdpb_inst_68_dout_w[15:0],sdpb_inst_68_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_68}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_196}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_68.READ_MODE = 1'b0;
defparam sdpb_inst_68.BIT_WIDTH_0 = 16;
defparam sdpb_inst_68.BIT_WIDTH_1 = 16;
defparam sdpb_inst_68.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_68.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_68.RESET_MODE = "SYNC";

SDPB sdpb_inst_69 (
    .DO({sdpb_inst_69_dout_w[15:0],sdpb_inst_69_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_69}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_197}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_69.READ_MODE = 1'b0;
defparam sdpb_inst_69.BIT_WIDTH_0 = 16;
defparam sdpb_inst_69.BIT_WIDTH_1 = 16;
defparam sdpb_inst_69.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_69.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_69.RESET_MODE = "SYNC";

SDPB sdpb_inst_70 (
    .DO({sdpb_inst_70_dout_w[15:0],sdpb_inst_70_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_70}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_198}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_70.READ_MODE = 1'b0;
defparam sdpb_inst_70.BIT_WIDTH_0 = 16;
defparam sdpb_inst_70.BIT_WIDTH_1 = 16;
defparam sdpb_inst_70.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_70.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_70.RESET_MODE = "SYNC";

SDPB sdpb_inst_71 (
    .DO({sdpb_inst_71_dout_w[15:0],sdpb_inst_71_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_71}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_199}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_71.READ_MODE = 1'b0;
defparam sdpb_inst_71.BIT_WIDTH_0 = 16;
defparam sdpb_inst_71.BIT_WIDTH_1 = 16;
defparam sdpb_inst_71.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_71.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_71.RESET_MODE = "SYNC";

SDPB sdpb_inst_72 (
    .DO({sdpb_inst_72_dout_w[15:0],sdpb_inst_72_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_72}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_200}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_72.READ_MODE = 1'b0;
defparam sdpb_inst_72.BIT_WIDTH_0 = 16;
defparam sdpb_inst_72.BIT_WIDTH_1 = 16;
defparam sdpb_inst_72.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_72.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_72.RESET_MODE = "SYNC";

SDPB sdpb_inst_73 (
    .DO({sdpb_inst_73_dout_w[15:0],sdpb_inst_73_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_73}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_201}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_73.READ_MODE = 1'b0;
defparam sdpb_inst_73.BIT_WIDTH_0 = 16;
defparam sdpb_inst_73.BIT_WIDTH_1 = 16;
defparam sdpb_inst_73.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_73.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_73.RESET_MODE = "SYNC";

SDPB sdpb_inst_74 (
    .DO({sdpb_inst_74_dout_w[15:0],sdpb_inst_74_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_74}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_202}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_74.READ_MODE = 1'b0;
defparam sdpb_inst_74.BIT_WIDTH_0 = 16;
defparam sdpb_inst_74.BIT_WIDTH_1 = 16;
defparam sdpb_inst_74.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_74.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_74.RESET_MODE = "SYNC";

SDPB sdpb_inst_75 (
    .DO({sdpb_inst_75_dout_w[15:0],sdpb_inst_75_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_75}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_203}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_75.READ_MODE = 1'b0;
defparam sdpb_inst_75.BIT_WIDTH_0 = 16;
defparam sdpb_inst_75.BIT_WIDTH_1 = 16;
defparam sdpb_inst_75.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_75.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_75.RESET_MODE = "SYNC";

SDPB sdpb_inst_76 (
    .DO({sdpb_inst_76_dout_w[15:0],sdpb_inst_76_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_76}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_204}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_76.READ_MODE = 1'b0;
defparam sdpb_inst_76.BIT_WIDTH_0 = 16;
defparam sdpb_inst_76.BIT_WIDTH_1 = 16;
defparam sdpb_inst_76.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_76.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_76.RESET_MODE = "SYNC";

SDPB sdpb_inst_77 (
    .DO({sdpb_inst_77_dout_w[15:0],sdpb_inst_77_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_77}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_205}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_77.READ_MODE = 1'b0;
defparam sdpb_inst_77.BIT_WIDTH_0 = 16;
defparam sdpb_inst_77.BIT_WIDTH_1 = 16;
defparam sdpb_inst_77.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_77.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_77.RESET_MODE = "SYNC";

SDPB sdpb_inst_78 (
    .DO({sdpb_inst_78_dout_w[15:0],sdpb_inst_78_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_78}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_206}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_78.READ_MODE = 1'b0;
defparam sdpb_inst_78.BIT_WIDTH_0 = 16;
defparam sdpb_inst_78.BIT_WIDTH_1 = 16;
defparam sdpb_inst_78.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_78.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_78.RESET_MODE = "SYNC";

SDPB sdpb_inst_79 (
    .DO({sdpb_inst_79_dout_w[15:0],sdpb_inst_79_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_79}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_207}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_79.READ_MODE = 1'b0;
defparam sdpb_inst_79.BIT_WIDTH_0 = 16;
defparam sdpb_inst_79.BIT_WIDTH_1 = 16;
defparam sdpb_inst_79.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_79.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_79.RESET_MODE = "SYNC";

SDPB sdpb_inst_80 (
    .DO({sdpb_inst_80_dout_w[15:0],sdpb_inst_80_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_80}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_208}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_80.READ_MODE = 1'b0;
defparam sdpb_inst_80.BIT_WIDTH_0 = 16;
defparam sdpb_inst_80.BIT_WIDTH_1 = 16;
defparam sdpb_inst_80.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_80.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_80.RESET_MODE = "SYNC";

SDPB sdpb_inst_81 (
    .DO({sdpb_inst_81_dout_w[15:0],sdpb_inst_81_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_81}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_209}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_81.READ_MODE = 1'b0;
defparam sdpb_inst_81.BIT_WIDTH_0 = 16;
defparam sdpb_inst_81.BIT_WIDTH_1 = 16;
defparam sdpb_inst_81.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_81.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_81.RESET_MODE = "SYNC";

SDPB sdpb_inst_82 (
    .DO({sdpb_inst_82_dout_w[15:0],sdpb_inst_82_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_82}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_210}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_82.READ_MODE = 1'b0;
defparam sdpb_inst_82.BIT_WIDTH_0 = 16;
defparam sdpb_inst_82.BIT_WIDTH_1 = 16;
defparam sdpb_inst_82.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_82.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_82.RESET_MODE = "SYNC";

SDPB sdpb_inst_83 (
    .DO({sdpb_inst_83_dout_w[15:0],sdpb_inst_83_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_83}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_211}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_83.READ_MODE = 1'b0;
defparam sdpb_inst_83.BIT_WIDTH_0 = 16;
defparam sdpb_inst_83.BIT_WIDTH_1 = 16;
defparam sdpb_inst_83.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_83.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_83.RESET_MODE = "SYNC";

SDPB sdpb_inst_84 (
    .DO({sdpb_inst_84_dout_w[15:0],sdpb_inst_84_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_84}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_212}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_84.READ_MODE = 1'b0;
defparam sdpb_inst_84.BIT_WIDTH_0 = 16;
defparam sdpb_inst_84.BIT_WIDTH_1 = 16;
defparam sdpb_inst_84.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_84.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_84.RESET_MODE = "SYNC";

SDPB sdpb_inst_85 (
    .DO({sdpb_inst_85_dout_w[15:0],sdpb_inst_85_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_85}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_213}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_85.READ_MODE = 1'b0;
defparam sdpb_inst_85.BIT_WIDTH_0 = 16;
defparam sdpb_inst_85.BIT_WIDTH_1 = 16;
defparam sdpb_inst_85.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_85.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_85.RESET_MODE = "SYNC";

SDPB sdpb_inst_86 (
    .DO({sdpb_inst_86_dout_w[15:0],sdpb_inst_86_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_86}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_214}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_86.READ_MODE = 1'b0;
defparam sdpb_inst_86.BIT_WIDTH_0 = 16;
defparam sdpb_inst_86.BIT_WIDTH_1 = 16;
defparam sdpb_inst_86.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_86.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_86.RESET_MODE = "SYNC";

SDPB sdpb_inst_87 (
    .DO({sdpb_inst_87_dout_w[15:0],sdpb_inst_87_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_87}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_215}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_87.READ_MODE = 1'b0;
defparam sdpb_inst_87.BIT_WIDTH_0 = 16;
defparam sdpb_inst_87.BIT_WIDTH_1 = 16;
defparam sdpb_inst_87.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_87.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_87.RESET_MODE = "SYNC";

SDPB sdpb_inst_88 (
    .DO({sdpb_inst_88_dout_w[15:0],sdpb_inst_88_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_88}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_216}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_88.READ_MODE = 1'b0;
defparam sdpb_inst_88.BIT_WIDTH_0 = 16;
defparam sdpb_inst_88.BIT_WIDTH_1 = 16;
defparam sdpb_inst_88.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_88.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_88.RESET_MODE = "SYNC";

SDPB sdpb_inst_89 (
    .DO({sdpb_inst_89_dout_w[15:0],sdpb_inst_89_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_89}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_217}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_89.READ_MODE = 1'b0;
defparam sdpb_inst_89.BIT_WIDTH_0 = 16;
defparam sdpb_inst_89.BIT_WIDTH_1 = 16;
defparam sdpb_inst_89.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_89.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_89.RESET_MODE = "SYNC";

SDPB sdpb_inst_90 (
    .DO({sdpb_inst_90_dout_w[15:0],sdpb_inst_90_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_90}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_218}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_90.READ_MODE = 1'b0;
defparam sdpb_inst_90.BIT_WIDTH_0 = 16;
defparam sdpb_inst_90.BIT_WIDTH_1 = 16;
defparam sdpb_inst_90.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_90.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_90.RESET_MODE = "SYNC";

SDPB sdpb_inst_91 (
    .DO({sdpb_inst_91_dout_w[15:0],sdpb_inst_91_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_91}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_219}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_91.READ_MODE = 1'b0;
defparam sdpb_inst_91.BIT_WIDTH_0 = 16;
defparam sdpb_inst_91.BIT_WIDTH_1 = 16;
defparam sdpb_inst_91.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_91.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_91.RESET_MODE = "SYNC";

SDPB sdpb_inst_92 (
    .DO({sdpb_inst_92_dout_w[15:0],sdpb_inst_92_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_92}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_220}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_92.READ_MODE = 1'b0;
defparam sdpb_inst_92.BIT_WIDTH_0 = 16;
defparam sdpb_inst_92.BIT_WIDTH_1 = 16;
defparam sdpb_inst_92.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_92.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_92.RESET_MODE = "SYNC";

SDPB sdpb_inst_93 (
    .DO({sdpb_inst_93_dout_w[15:0],sdpb_inst_93_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_93}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_221}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_93.READ_MODE = 1'b0;
defparam sdpb_inst_93.BIT_WIDTH_0 = 16;
defparam sdpb_inst_93.BIT_WIDTH_1 = 16;
defparam sdpb_inst_93.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_93.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_93.RESET_MODE = "SYNC";

SDPB sdpb_inst_94 (
    .DO({sdpb_inst_94_dout_w[15:0],sdpb_inst_94_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_94}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_222}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_94.READ_MODE = 1'b0;
defparam sdpb_inst_94.BIT_WIDTH_0 = 16;
defparam sdpb_inst_94.BIT_WIDTH_1 = 16;
defparam sdpb_inst_94.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_94.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_94.RESET_MODE = "SYNC";

SDPB sdpb_inst_95 (
    .DO({sdpb_inst_95_dout_w[15:0],sdpb_inst_95_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_95}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_223}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_95.READ_MODE = 1'b0;
defparam sdpb_inst_95.BIT_WIDTH_0 = 16;
defparam sdpb_inst_95.BIT_WIDTH_1 = 16;
defparam sdpb_inst_95.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_95.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_95.RESET_MODE = "SYNC";

SDPB sdpb_inst_96 (
    .DO({sdpb_inst_96_dout_w[15:0],sdpb_inst_96_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_96}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_224}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_96.READ_MODE = 1'b0;
defparam sdpb_inst_96.BIT_WIDTH_0 = 16;
defparam sdpb_inst_96.BIT_WIDTH_1 = 16;
defparam sdpb_inst_96.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_96.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_96.RESET_MODE = "SYNC";

SDPB sdpb_inst_97 (
    .DO({sdpb_inst_97_dout_w[15:0],sdpb_inst_97_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_97}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_225}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_97.READ_MODE = 1'b0;
defparam sdpb_inst_97.BIT_WIDTH_0 = 16;
defparam sdpb_inst_97.BIT_WIDTH_1 = 16;
defparam sdpb_inst_97.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_97.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_97.RESET_MODE = "SYNC";

SDPB sdpb_inst_98 (
    .DO({sdpb_inst_98_dout_w[15:0],sdpb_inst_98_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_98}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_226}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_98.READ_MODE = 1'b0;
defparam sdpb_inst_98.BIT_WIDTH_0 = 16;
defparam sdpb_inst_98.BIT_WIDTH_1 = 16;
defparam sdpb_inst_98.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_98.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_98.RESET_MODE = "SYNC";

SDPB sdpb_inst_99 (
    .DO({sdpb_inst_99_dout_w[15:0],sdpb_inst_99_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_99}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_227}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_99.READ_MODE = 1'b0;
defparam sdpb_inst_99.BIT_WIDTH_0 = 16;
defparam sdpb_inst_99.BIT_WIDTH_1 = 16;
defparam sdpb_inst_99.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_99.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_99.RESET_MODE = "SYNC";

SDPB sdpb_inst_100 (
    .DO({sdpb_inst_100_dout_w[15:0],sdpb_inst_100_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_100}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_228}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_100.READ_MODE = 1'b0;
defparam sdpb_inst_100.BIT_WIDTH_0 = 16;
defparam sdpb_inst_100.BIT_WIDTH_1 = 16;
defparam sdpb_inst_100.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_100.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_100.RESET_MODE = "SYNC";

SDPB sdpb_inst_101 (
    .DO({sdpb_inst_101_dout_w[15:0],sdpb_inst_101_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_101}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_229}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_101.READ_MODE = 1'b0;
defparam sdpb_inst_101.BIT_WIDTH_0 = 16;
defparam sdpb_inst_101.BIT_WIDTH_1 = 16;
defparam sdpb_inst_101.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_101.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_101.RESET_MODE = "SYNC";

SDPB sdpb_inst_102 (
    .DO({sdpb_inst_102_dout_w[15:0],sdpb_inst_102_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_102}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_230}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_102.READ_MODE = 1'b0;
defparam sdpb_inst_102.BIT_WIDTH_0 = 16;
defparam sdpb_inst_102.BIT_WIDTH_1 = 16;
defparam sdpb_inst_102.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_102.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_102.RESET_MODE = "SYNC";

SDPB sdpb_inst_103 (
    .DO({sdpb_inst_103_dout_w[15:0],sdpb_inst_103_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_103}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_231}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_103.READ_MODE = 1'b0;
defparam sdpb_inst_103.BIT_WIDTH_0 = 16;
defparam sdpb_inst_103.BIT_WIDTH_1 = 16;
defparam sdpb_inst_103.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_103.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_103.RESET_MODE = "SYNC";

SDPB sdpb_inst_104 (
    .DO({sdpb_inst_104_dout_w[15:0],sdpb_inst_104_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_104}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_232}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_104.READ_MODE = 1'b0;
defparam sdpb_inst_104.BIT_WIDTH_0 = 16;
defparam sdpb_inst_104.BIT_WIDTH_1 = 16;
defparam sdpb_inst_104.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_104.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_104.RESET_MODE = "SYNC";

SDPB sdpb_inst_105 (
    .DO({sdpb_inst_105_dout_w[15:0],sdpb_inst_105_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_105}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_233}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_105.READ_MODE = 1'b0;
defparam sdpb_inst_105.BIT_WIDTH_0 = 16;
defparam sdpb_inst_105.BIT_WIDTH_1 = 16;
defparam sdpb_inst_105.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_105.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_105.RESET_MODE = "SYNC";

SDPB sdpb_inst_106 (
    .DO({sdpb_inst_106_dout_w[15:0],sdpb_inst_106_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_106}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_234}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_106.READ_MODE = 1'b0;
defparam sdpb_inst_106.BIT_WIDTH_0 = 16;
defparam sdpb_inst_106.BIT_WIDTH_1 = 16;
defparam sdpb_inst_106.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_106.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_106.RESET_MODE = "SYNC";

SDPB sdpb_inst_107 (
    .DO({sdpb_inst_107_dout_w[15:0],sdpb_inst_107_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_107}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_235}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_107.READ_MODE = 1'b0;
defparam sdpb_inst_107.BIT_WIDTH_0 = 16;
defparam sdpb_inst_107.BIT_WIDTH_1 = 16;
defparam sdpb_inst_107.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_107.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_107.RESET_MODE = "SYNC";

SDPB sdpb_inst_108 (
    .DO({sdpb_inst_108_dout_w[15:0],sdpb_inst_108_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_108}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_236}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_108.READ_MODE = 1'b0;
defparam sdpb_inst_108.BIT_WIDTH_0 = 16;
defparam sdpb_inst_108.BIT_WIDTH_1 = 16;
defparam sdpb_inst_108.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_108.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_108.RESET_MODE = "SYNC";

SDPB sdpb_inst_109 (
    .DO({sdpb_inst_109_dout_w[15:0],sdpb_inst_109_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_109}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_237}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_109.READ_MODE = 1'b0;
defparam sdpb_inst_109.BIT_WIDTH_0 = 16;
defparam sdpb_inst_109.BIT_WIDTH_1 = 16;
defparam sdpb_inst_109.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_109.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_109.RESET_MODE = "SYNC";

SDPB sdpb_inst_110 (
    .DO({sdpb_inst_110_dout_w[15:0],sdpb_inst_110_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_110}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_238}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_110.READ_MODE = 1'b0;
defparam sdpb_inst_110.BIT_WIDTH_0 = 16;
defparam sdpb_inst_110.BIT_WIDTH_1 = 16;
defparam sdpb_inst_110.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_110.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_110.RESET_MODE = "SYNC";

SDPB sdpb_inst_111 (
    .DO({sdpb_inst_111_dout_w[15:0],sdpb_inst_111_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_111}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_239}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_111.READ_MODE = 1'b0;
defparam sdpb_inst_111.BIT_WIDTH_0 = 16;
defparam sdpb_inst_111.BIT_WIDTH_1 = 16;
defparam sdpb_inst_111.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_111.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_111.RESET_MODE = "SYNC";

SDPB sdpb_inst_112 (
    .DO({sdpb_inst_112_dout_w[15:0],sdpb_inst_112_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_112}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_240}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_112.READ_MODE = 1'b0;
defparam sdpb_inst_112.BIT_WIDTH_0 = 16;
defparam sdpb_inst_112.BIT_WIDTH_1 = 16;
defparam sdpb_inst_112.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_112.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_112.RESET_MODE = "SYNC";

SDPB sdpb_inst_113 (
    .DO({sdpb_inst_113_dout_w[15:0],sdpb_inst_113_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_113}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_241}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_113.READ_MODE = 1'b0;
defparam sdpb_inst_113.BIT_WIDTH_0 = 16;
defparam sdpb_inst_113.BIT_WIDTH_1 = 16;
defparam sdpb_inst_113.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_113.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_113.RESET_MODE = "SYNC";

SDPB sdpb_inst_114 (
    .DO({sdpb_inst_114_dout_w[15:0],sdpb_inst_114_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_114}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_242}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_114.READ_MODE = 1'b0;
defparam sdpb_inst_114.BIT_WIDTH_0 = 16;
defparam sdpb_inst_114.BIT_WIDTH_1 = 16;
defparam sdpb_inst_114.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_114.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_114.RESET_MODE = "SYNC";

SDPB sdpb_inst_115 (
    .DO({sdpb_inst_115_dout_w[15:0],sdpb_inst_115_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_115}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_243}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_115.READ_MODE = 1'b0;
defparam sdpb_inst_115.BIT_WIDTH_0 = 16;
defparam sdpb_inst_115.BIT_WIDTH_1 = 16;
defparam sdpb_inst_115.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_115.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_115.RESET_MODE = "SYNC";

SDPB sdpb_inst_116 (
    .DO({sdpb_inst_116_dout_w[15:0],sdpb_inst_116_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_116}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_244}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_116.READ_MODE = 1'b0;
defparam sdpb_inst_116.BIT_WIDTH_0 = 16;
defparam sdpb_inst_116.BIT_WIDTH_1 = 16;
defparam sdpb_inst_116.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_116.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_116.RESET_MODE = "SYNC";

SDPB sdpb_inst_117 (
    .DO({sdpb_inst_117_dout_w[15:0],sdpb_inst_117_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_117}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_245}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_117.READ_MODE = 1'b0;
defparam sdpb_inst_117.BIT_WIDTH_0 = 16;
defparam sdpb_inst_117.BIT_WIDTH_1 = 16;
defparam sdpb_inst_117.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_117.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_117.RESET_MODE = "SYNC";

SDPB sdpb_inst_118 (
    .DO({sdpb_inst_118_dout_w[15:0],sdpb_inst_118_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_118}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_246}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_118.READ_MODE = 1'b0;
defparam sdpb_inst_118.BIT_WIDTH_0 = 16;
defparam sdpb_inst_118.BIT_WIDTH_1 = 16;
defparam sdpb_inst_118.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_118.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_118.RESET_MODE = "SYNC";

SDPB sdpb_inst_119 (
    .DO({sdpb_inst_119_dout_w[15:0],sdpb_inst_119_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_119}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_247}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_119.READ_MODE = 1'b0;
defparam sdpb_inst_119.BIT_WIDTH_0 = 16;
defparam sdpb_inst_119.BIT_WIDTH_1 = 16;
defparam sdpb_inst_119.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_119.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_119.RESET_MODE = "SYNC";

SDPB sdpb_inst_120 (
    .DO({sdpb_inst_120_dout_w[15:0],sdpb_inst_120_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_120}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_248}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_120.READ_MODE = 1'b0;
defparam sdpb_inst_120.BIT_WIDTH_0 = 16;
defparam sdpb_inst_120.BIT_WIDTH_1 = 16;
defparam sdpb_inst_120.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_120.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_120.RESET_MODE = "SYNC";

SDPB sdpb_inst_121 (
    .DO({sdpb_inst_121_dout_w[15:0],sdpb_inst_121_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_121}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_249}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_121.READ_MODE = 1'b0;
defparam sdpb_inst_121.BIT_WIDTH_0 = 16;
defparam sdpb_inst_121.BIT_WIDTH_1 = 16;
defparam sdpb_inst_121.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_121.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_121.RESET_MODE = "SYNC";

SDPB sdpb_inst_122 (
    .DO({sdpb_inst_122_dout_w[15:0],sdpb_inst_122_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_122}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_250}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_122.READ_MODE = 1'b0;
defparam sdpb_inst_122.BIT_WIDTH_0 = 16;
defparam sdpb_inst_122.BIT_WIDTH_1 = 16;
defparam sdpb_inst_122.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_122.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_122.RESET_MODE = "SYNC";

SDPB sdpb_inst_123 (
    .DO({sdpb_inst_123_dout_w[15:0],sdpb_inst_123_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_123}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_251}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_123.READ_MODE = 1'b0;
defparam sdpb_inst_123.BIT_WIDTH_0 = 16;
defparam sdpb_inst_123.BIT_WIDTH_1 = 16;
defparam sdpb_inst_123.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_123.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_123.RESET_MODE = "SYNC";

SDPB sdpb_inst_124 (
    .DO({sdpb_inst_124_dout_w[15:0],sdpb_inst_124_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_124}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_252}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_124.READ_MODE = 1'b0;
defparam sdpb_inst_124.BIT_WIDTH_0 = 16;
defparam sdpb_inst_124.BIT_WIDTH_1 = 16;
defparam sdpb_inst_124.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_124.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_124.RESET_MODE = "SYNC";

SDPB sdpb_inst_125 (
    .DO({sdpb_inst_125_dout_w[15:0],sdpb_inst_125_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_125}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_253}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_125.READ_MODE = 1'b0;
defparam sdpb_inst_125.BIT_WIDTH_0 = 16;
defparam sdpb_inst_125.BIT_WIDTH_1 = 16;
defparam sdpb_inst_125.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_125.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_125.RESET_MODE = "SYNC";

SDPB sdpb_inst_126 (
    .DO({sdpb_inst_126_dout_w[15:0],sdpb_inst_126_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_126}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_254}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_126.READ_MODE = 1'b0;
defparam sdpb_inst_126.BIT_WIDTH_0 = 16;
defparam sdpb_inst_126.BIT_WIDTH_1 = 16;
defparam sdpb_inst_126.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_126.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_126.RESET_MODE = "SYNC";

SDPB sdpb_inst_127 (
    .DO({sdpb_inst_127_dout_w[15:0],sdpb_inst_127_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_127}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_255}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_127.READ_MODE = 1'b0;
defparam sdpb_inst_127.BIT_WIDTH_0 = 16;
defparam sdpb_inst_127.BIT_WIDTH_1 = 16;
defparam sdpb_inst_127.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_127.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_127.RESET_MODE = "SYNC";

SDPB sdpb_inst_128 (
    .DO({sdpb_inst_128_dout_w[15:0],sdpb_inst_128_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_128}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_128.READ_MODE = 1'b0;
defparam sdpb_inst_128.BIT_WIDTH_0 = 16;
defparam sdpb_inst_128.BIT_WIDTH_1 = 16;
defparam sdpb_inst_128.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_128.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_128.RESET_MODE = "SYNC";

SDPB sdpb_inst_129 (
    .DO({sdpb_inst_129_dout_w[15:0],sdpb_inst_129_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_129}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_129.READ_MODE = 1'b0;
defparam sdpb_inst_129.BIT_WIDTH_0 = 16;
defparam sdpb_inst_129.BIT_WIDTH_1 = 16;
defparam sdpb_inst_129.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_129.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_129.RESET_MODE = "SYNC";

SDPB sdpb_inst_130 (
    .DO({sdpb_inst_130_dout_w[15:0],sdpb_inst_130_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_130}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_130.READ_MODE = 1'b0;
defparam sdpb_inst_130.BIT_WIDTH_0 = 16;
defparam sdpb_inst_130.BIT_WIDTH_1 = 16;
defparam sdpb_inst_130.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_130.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_130.RESET_MODE = "SYNC";

SDPB sdpb_inst_131 (
    .DO({sdpb_inst_131_dout_w[15:0],sdpb_inst_131_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_131}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_131.READ_MODE = 1'b0;
defparam sdpb_inst_131.BIT_WIDTH_0 = 16;
defparam sdpb_inst_131.BIT_WIDTH_1 = 16;
defparam sdpb_inst_131.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_131.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_131.RESET_MODE = "SYNC";

SDPB sdpb_inst_132 (
    .DO({sdpb_inst_132_dout_w[15:0],sdpb_inst_132_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_132}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_132.READ_MODE = 1'b0;
defparam sdpb_inst_132.BIT_WIDTH_0 = 16;
defparam sdpb_inst_132.BIT_WIDTH_1 = 16;
defparam sdpb_inst_132.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_132.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_132.RESET_MODE = "SYNC";

SDPB sdpb_inst_133 (
    .DO({sdpb_inst_133_dout_w[15:0],sdpb_inst_133_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_133}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_133.READ_MODE = 1'b0;
defparam sdpb_inst_133.BIT_WIDTH_0 = 16;
defparam sdpb_inst_133.BIT_WIDTH_1 = 16;
defparam sdpb_inst_133.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_133.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_133.RESET_MODE = "SYNC";

SDPB sdpb_inst_134 (
    .DO({sdpb_inst_134_dout_w[15:0],sdpb_inst_134_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_134}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_134.READ_MODE = 1'b0;
defparam sdpb_inst_134.BIT_WIDTH_0 = 16;
defparam sdpb_inst_134.BIT_WIDTH_1 = 16;
defparam sdpb_inst_134.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_134.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_134.RESET_MODE = "SYNC";

SDPB sdpb_inst_135 (
    .DO({sdpb_inst_135_dout_w[15:0],sdpb_inst_135_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_135}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_135.READ_MODE = 1'b0;
defparam sdpb_inst_135.BIT_WIDTH_0 = 16;
defparam sdpb_inst_135.BIT_WIDTH_1 = 16;
defparam sdpb_inst_135.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_135.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_135.RESET_MODE = "SYNC";

SDPB sdpb_inst_136 (
    .DO({sdpb_inst_136_dout_w[15:0],sdpb_inst_136_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_136}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_136.READ_MODE = 1'b0;
defparam sdpb_inst_136.BIT_WIDTH_0 = 16;
defparam sdpb_inst_136.BIT_WIDTH_1 = 16;
defparam sdpb_inst_136.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_136.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_136.RESET_MODE = "SYNC";

SDPB sdpb_inst_137 (
    .DO({sdpb_inst_137_dout_w[15:0],sdpb_inst_137_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_137}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_137.READ_MODE = 1'b0;
defparam sdpb_inst_137.BIT_WIDTH_0 = 16;
defparam sdpb_inst_137.BIT_WIDTH_1 = 16;
defparam sdpb_inst_137.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_137.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_137.RESET_MODE = "SYNC";

SDPB sdpb_inst_138 (
    .DO({sdpb_inst_138_dout_w[15:0],sdpb_inst_138_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_138}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_138.READ_MODE = 1'b0;
defparam sdpb_inst_138.BIT_WIDTH_0 = 16;
defparam sdpb_inst_138.BIT_WIDTH_1 = 16;
defparam sdpb_inst_138.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_138.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_138.RESET_MODE = "SYNC";

SDPB sdpb_inst_139 (
    .DO({sdpb_inst_139_dout_w[15:0],sdpb_inst_139_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_139}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_139.READ_MODE = 1'b0;
defparam sdpb_inst_139.BIT_WIDTH_0 = 16;
defparam sdpb_inst_139.BIT_WIDTH_1 = 16;
defparam sdpb_inst_139.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_139.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_139.RESET_MODE = "SYNC";

SDPB sdpb_inst_140 (
    .DO({sdpb_inst_140_dout_w[15:0],sdpb_inst_140_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_140}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_140.READ_MODE = 1'b0;
defparam sdpb_inst_140.BIT_WIDTH_0 = 16;
defparam sdpb_inst_140.BIT_WIDTH_1 = 16;
defparam sdpb_inst_140.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_140.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_140.RESET_MODE = "SYNC";

SDPB sdpb_inst_141 (
    .DO({sdpb_inst_141_dout_w[15:0],sdpb_inst_141_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_141}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_141.READ_MODE = 1'b0;
defparam sdpb_inst_141.BIT_WIDTH_0 = 16;
defparam sdpb_inst_141.BIT_WIDTH_1 = 16;
defparam sdpb_inst_141.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_141.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_141.RESET_MODE = "SYNC";

SDPB sdpb_inst_142 (
    .DO({sdpb_inst_142_dout_w[15:0],sdpb_inst_142_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_142}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_142.READ_MODE = 1'b0;
defparam sdpb_inst_142.BIT_WIDTH_0 = 16;
defparam sdpb_inst_142.BIT_WIDTH_1 = 16;
defparam sdpb_inst_142.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_142.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_142.RESET_MODE = "SYNC";

SDPB sdpb_inst_143 (
    .DO({sdpb_inst_143_dout_w[15:0],sdpb_inst_143_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_143}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_143.READ_MODE = 1'b0;
defparam sdpb_inst_143.BIT_WIDTH_0 = 16;
defparam sdpb_inst_143.BIT_WIDTH_1 = 16;
defparam sdpb_inst_143.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_143.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_143.RESET_MODE = "SYNC";

SDPB sdpb_inst_144 (
    .DO({sdpb_inst_144_dout_w[15:0],sdpb_inst_144_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_16}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_144}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_144.READ_MODE = 1'b0;
defparam sdpb_inst_144.BIT_WIDTH_0 = 16;
defparam sdpb_inst_144.BIT_WIDTH_1 = 16;
defparam sdpb_inst_144.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_144.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_144.RESET_MODE = "SYNC";

SDPB sdpb_inst_145 (
    .DO({sdpb_inst_145_dout_w[15:0],sdpb_inst_145_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_17}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_145}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_145.READ_MODE = 1'b0;
defparam sdpb_inst_145.BIT_WIDTH_0 = 16;
defparam sdpb_inst_145.BIT_WIDTH_1 = 16;
defparam sdpb_inst_145.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_145.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_145.RESET_MODE = "SYNC";

SDPB sdpb_inst_146 (
    .DO({sdpb_inst_146_dout_w[15:0],sdpb_inst_146_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_18}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_146}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_146.READ_MODE = 1'b0;
defparam sdpb_inst_146.BIT_WIDTH_0 = 16;
defparam sdpb_inst_146.BIT_WIDTH_1 = 16;
defparam sdpb_inst_146.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_146.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_146.RESET_MODE = "SYNC";

SDPB sdpb_inst_147 (
    .DO({sdpb_inst_147_dout_w[15:0],sdpb_inst_147_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_19}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_147}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_147.READ_MODE = 1'b0;
defparam sdpb_inst_147.BIT_WIDTH_0 = 16;
defparam sdpb_inst_147.BIT_WIDTH_1 = 16;
defparam sdpb_inst_147.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_147.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_147.RESET_MODE = "SYNC";

SDPB sdpb_inst_148 (
    .DO({sdpb_inst_148_dout_w[15:0],sdpb_inst_148_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_20}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_148}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_148.READ_MODE = 1'b0;
defparam sdpb_inst_148.BIT_WIDTH_0 = 16;
defparam sdpb_inst_148.BIT_WIDTH_1 = 16;
defparam sdpb_inst_148.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_148.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_148.RESET_MODE = "SYNC";

SDPB sdpb_inst_149 (
    .DO({sdpb_inst_149_dout_w[15:0],sdpb_inst_149_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_21}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_149}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_149.READ_MODE = 1'b0;
defparam sdpb_inst_149.BIT_WIDTH_0 = 16;
defparam sdpb_inst_149.BIT_WIDTH_1 = 16;
defparam sdpb_inst_149.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_149.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_149.RESET_MODE = "SYNC";

SDPB sdpb_inst_150 (
    .DO({sdpb_inst_150_dout_w[15:0],sdpb_inst_150_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_22}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_150}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_150.READ_MODE = 1'b0;
defparam sdpb_inst_150.BIT_WIDTH_0 = 16;
defparam sdpb_inst_150.BIT_WIDTH_1 = 16;
defparam sdpb_inst_150.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_150.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_150.RESET_MODE = "SYNC";

SDPB sdpb_inst_151 (
    .DO({sdpb_inst_151_dout_w[15:0],sdpb_inst_151_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_23}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_151}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_151.READ_MODE = 1'b0;
defparam sdpb_inst_151.BIT_WIDTH_0 = 16;
defparam sdpb_inst_151.BIT_WIDTH_1 = 16;
defparam sdpb_inst_151.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_151.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_151.RESET_MODE = "SYNC";

SDPB sdpb_inst_152 (
    .DO({sdpb_inst_152_dout_w[15:0],sdpb_inst_152_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_24}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_152}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_152.READ_MODE = 1'b0;
defparam sdpb_inst_152.BIT_WIDTH_0 = 16;
defparam sdpb_inst_152.BIT_WIDTH_1 = 16;
defparam sdpb_inst_152.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_152.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_152.RESET_MODE = "SYNC";

SDPB sdpb_inst_153 (
    .DO({sdpb_inst_153_dout_w[15:0],sdpb_inst_153_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_25}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_153}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_153.READ_MODE = 1'b0;
defparam sdpb_inst_153.BIT_WIDTH_0 = 16;
defparam sdpb_inst_153.BIT_WIDTH_1 = 16;
defparam sdpb_inst_153.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_153.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_153.RESET_MODE = "SYNC";

SDPB sdpb_inst_154 (
    .DO({sdpb_inst_154_dout_w[15:0],sdpb_inst_154_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_26}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_154}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_154.READ_MODE = 1'b0;
defparam sdpb_inst_154.BIT_WIDTH_0 = 16;
defparam sdpb_inst_154.BIT_WIDTH_1 = 16;
defparam sdpb_inst_154.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_154.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_154.RESET_MODE = "SYNC";

SDPB sdpb_inst_155 (
    .DO({sdpb_inst_155_dout_w[15:0],sdpb_inst_155_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_27}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_155}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_155.READ_MODE = 1'b0;
defparam sdpb_inst_155.BIT_WIDTH_0 = 16;
defparam sdpb_inst_155.BIT_WIDTH_1 = 16;
defparam sdpb_inst_155.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_155.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_155.RESET_MODE = "SYNC";

SDPB sdpb_inst_156 (
    .DO({sdpb_inst_156_dout_w[15:0],sdpb_inst_156_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_28}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_156}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_156.READ_MODE = 1'b0;
defparam sdpb_inst_156.BIT_WIDTH_0 = 16;
defparam sdpb_inst_156.BIT_WIDTH_1 = 16;
defparam sdpb_inst_156.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_156.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_156.RESET_MODE = "SYNC";

SDPB sdpb_inst_157 (
    .DO({sdpb_inst_157_dout_w[15:0],sdpb_inst_157_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_29}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_157}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_157.READ_MODE = 1'b0;
defparam sdpb_inst_157.BIT_WIDTH_0 = 16;
defparam sdpb_inst_157.BIT_WIDTH_1 = 16;
defparam sdpb_inst_157.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_157.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_157.RESET_MODE = "SYNC";

SDPB sdpb_inst_158 (
    .DO({sdpb_inst_158_dout_w[15:0],sdpb_inst_158_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_30}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_158}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_158.READ_MODE = 1'b0;
defparam sdpb_inst_158.BIT_WIDTH_0 = 16;
defparam sdpb_inst_158.BIT_WIDTH_1 = 16;
defparam sdpb_inst_158.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_158.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_158.RESET_MODE = "SYNC";

SDPB sdpb_inst_159 (
    .DO({sdpb_inst_159_dout_w[15:0],sdpb_inst_159_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_31}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_159}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_159.READ_MODE = 1'b0;
defparam sdpb_inst_159.BIT_WIDTH_0 = 16;
defparam sdpb_inst_159.BIT_WIDTH_1 = 16;
defparam sdpb_inst_159.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_159.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_159.RESET_MODE = "SYNC";

SDPB sdpb_inst_160 (
    .DO({sdpb_inst_160_dout_w[15:0],sdpb_inst_160_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_32}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_160}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_160.READ_MODE = 1'b0;
defparam sdpb_inst_160.BIT_WIDTH_0 = 16;
defparam sdpb_inst_160.BIT_WIDTH_1 = 16;
defparam sdpb_inst_160.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_160.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_160.RESET_MODE = "SYNC";

SDPB sdpb_inst_161 (
    .DO({sdpb_inst_161_dout_w[15:0],sdpb_inst_161_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_33}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_161}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_161.READ_MODE = 1'b0;
defparam sdpb_inst_161.BIT_WIDTH_0 = 16;
defparam sdpb_inst_161.BIT_WIDTH_1 = 16;
defparam sdpb_inst_161.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_161.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_161.RESET_MODE = "SYNC";

SDPB sdpb_inst_162 (
    .DO({sdpb_inst_162_dout_w[15:0],sdpb_inst_162_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_34}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_162}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_162.READ_MODE = 1'b0;
defparam sdpb_inst_162.BIT_WIDTH_0 = 16;
defparam sdpb_inst_162.BIT_WIDTH_1 = 16;
defparam sdpb_inst_162.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_162.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_162.RESET_MODE = "SYNC";

SDPB sdpb_inst_163 (
    .DO({sdpb_inst_163_dout_w[15:0],sdpb_inst_163_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_35}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_163}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_163.READ_MODE = 1'b0;
defparam sdpb_inst_163.BIT_WIDTH_0 = 16;
defparam sdpb_inst_163.BIT_WIDTH_1 = 16;
defparam sdpb_inst_163.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_163.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_163.RESET_MODE = "SYNC";

SDPB sdpb_inst_164 (
    .DO({sdpb_inst_164_dout_w[15:0],sdpb_inst_164_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_36}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_164}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_164.READ_MODE = 1'b0;
defparam sdpb_inst_164.BIT_WIDTH_0 = 16;
defparam sdpb_inst_164.BIT_WIDTH_1 = 16;
defparam sdpb_inst_164.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_164.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_164.RESET_MODE = "SYNC";

SDPB sdpb_inst_165 (
    .DO({sdpb_inst_165_dout_w[15:0],sdpb_inst_165_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_37}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_165}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_165.READ_MODE = 1'b0;
defparam sdpb_inst_165.BIT_WIDTH_0 = 16;
defparam sdpb_inst_165.BIT_WIDTH_1 = 16;
defparam sdpb_inst_165.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_165.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_165.RESET_MODE = "SYNC";

SDPB sdpb_inst_166 (
    .DO({sdpb_inst_166_dout_w[15:0],sdpb_inst_166_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_38}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_166}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_166.READ_MODE = 1'b0;
defparam sdpb_inst_166.BIT_WIDTH_0 = 16;
defparam sdpb_inst_166.BIT_WIDTH_1 = 16;
defparam sdpb_inst_166.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_166.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_166.RESET_MODE = "SYNC";

SDPB sdpb_inst_167 (
    .DO({sdpb_inst_167_dout_w[15:0],sdpb_inst_167_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_39}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_167}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_167.READ_MODE = 1'b0;
defparam sdpb_inst_167.BIT_WIDTH_0 = 16;
defparam sdpb_inst_167.BIT_WIDTH_1 = 16;
defparam sdpb_inst_167.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_167.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_167.RESET_MODE = "SYNC";

SDPB sdpb_inst_168 (
    .DO({sdpb_inst_168_dout_w[15:0],sdpb_inst_168_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_40}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_168}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_168.READ_MODE = 1'b0;
defparam sdpb_inst_168.BIT_WIDTH_0 = 16;
defparam sdpb_inst_168.BIT_WIDTH_1 = 16;
defparam sdpb_inst_168.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_168.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_168.RESET_MODE = "SYNC";

SDPB sdpb_inst_169 (
    .DO({sdpb_inst_169_dout_w[15:0],sdpb_inst_169_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_41}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_169}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_169.READ_MODE = 1'b0;
defparam sdpb_inst_169.BIT_WIDTH_0 = 16;
defparam sdpb_inst_169.BIT_WIDTH_1 = 16;
defparam sdpb_inst_169.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_169.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_169.RESET_MODE = "SYNC";

SDPB sdpb_inst_170 (
    .DO({sdpb_inst_170_dout_w[15:0],sdpb_inst_170_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_42}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_170}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_170.READ_MODE = 1'b0;
defparam sdpb_inst_170.BIT_WIDTH_0 = 16;
defparam sdpb_inst_170.BIT_WIDTH_1 = 16;
defparam sdpb_inst_170.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_170.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_170.RESET_MODE = "SYNC";

SDPB sdpb_inst_171 (
    .DO({sdpb_inst_171_dout_w[15:0],sdpb_inst_171_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_43}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_171}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_171.READ_MODE = 1'b0;
defparam sdpb_inst_171.BIT_WIDTH_0 = 16;
defparam sdpb_inst_171.BIT_WIDTH_1 = 16;
defparam sdpb_inst_171.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_171.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_171.RESET_MODE = "SYNC";

SDPB sdpb_inst_172 (
    .DO({sdpb_inst_172_dout_w[15:0],sdpb_inst_172_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_44}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_172}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_172.READ_MODE = 1'b0;
defparam sdpb_inst_172.BIT_WIDTH_0 = 16;
defparam sdpb_inst_172.BIT_WIDTH_1 = 16;
defparam sdpb_inst_172.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_172.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_172.RESET_MODE = "SYNC";

SDPB sdpb_inst_173 (
    .DO({sdpb_inst_173_dout_w[15:0],sdpb_inst_173_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_45}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_173}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_173.READ_MODE = 1'b0;
defparam sdpb_inst_173.BIT_WIDTH_0 = 16;
defparam sdpb_inst_173.BIT_WIDTH_1 = 16;
defparam sdpb_inst_173.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_173.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_173.RESET_MODE = "SYNC";

SDPB sdpb_inst_174 (
    .DO({sdpb_inst_174_dout_w[15:0],sdpb_inst_174_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_46}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_174}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_174.READ_MODE = 1'b0;
defparam sdpb_inst_174.BIT_WIDTH_0 = 16;
defparam sdpb_inst_174.BIT_WIDTH_1 = 16;
defparam sdpb_inst_174.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_174.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_174.RESET_MODE = "SYNC";

SDPB sdpb_inst_175 (
    .DO({sdpb_inst_175_dout_w[15:0],sdpb_inst_175_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_47}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_175}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_175.READ_MODE = 1'b0;
defparam sdpb_inst_175.BIT_WIDTH_0 = 16;
defparam sdpb_inst_175.BIT_WIDTH_1 = 16;
defparam sdpb_inst_175.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_175.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_175.RESET_MODE = "SYNC";

SDPB sdpb_inst_176 (
    .DO({sdpb_inst_176_dout_w[15:0],sdpb_inst_176_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_48}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_176}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_176.READ_MODE = 1'b0;
defparam sdpb_inst_176.BIT_WIDTH_0 = 16;
defparam sdpb_inst_176.BIT_WIDTH_1 = 16;
defparam sdpb_inst_176.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_176.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_176.RESET_MODE = "SYNC";

SDPB sdpb_inst_177 (
    .DO({sdpb_inst_177_dout_w[15:0],sdpb_inst_177_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_49}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_177}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_177.READ_MODE = 1'b0;
defparam sdpb_inst_177.BIT_WIDTH_0 = 16;
defparam sdpb_inst_177.BIT_WIDTH_1 = 16;
defparam sdpb_inst_177.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_177.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_177.RESET_MODE = "SYNC";

SDPB sdpb_inst_178 (
    .DO({sdpb_inst_178_dout_w[15:0],sdpb_inst_178_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_50}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_178}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_178.READ_MODE = 1'b0;
defparam sdpb_inst_178.BIT_WIDTH_0 = 16;
defparam sdpb_inst_178.BIT_WIDTH_1 = 16;
defparam sdpb_inst_178.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_178.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_178.RESET_MODE = "SYNC";

SDPB sdpb_inst_179 (
    .DO({sdpb_inst_179_dout_w[15:0],sdpb_inst_179_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_51}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_179}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_179.READ_MODE = 1'b0;
defparam sdpb_inst_179.BIT_WIDTH_0 = 16;
defparam sdpb_inst_179.BIT_WIDTH_1 = 16;
defparam sdpb_inst_179.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_179.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_179.RESET_MODE = "SYNC";

SDPB sdpb_inst_180 (
    .DO({sdpb_inst_180_dout_w[15:0],sdpb_inst_180_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_52}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_180}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_180.READ_MODE = 1'b0;
defparam sdpb_inst_180.BIT_WIDTH_0 = 16;
defparam sdpb_inst_180.BIT_WIDTH_1 = 16;
defparam sdpb_inst_180.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_180.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_180.RESET_MODE = "SYNC";

SDPB sdpb_inst_181 (
    .DO({sdpb_inst_181_dout_w[15:0],sdpb_inst_181_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_53}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_181}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_181.READ_MODE = 1'b0;
defparam sdpb_inst_181.BIT_WIDTH_0 = 16;
defparam sdpb_inst_181.BIT_WIDTH_1 = 16;
defparam sdpb_inst_181.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_181.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_181.RESET_MODE = "SYNC";

SDPB sdpb_inst_182 (
    .DO({sdpb_inst_182_dout_w[15:0],sdpb_inst_182_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_54}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_182}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_182.READ_MODE = 1'b0;
defparam sdpb_inst_182.BIT_WIDTH_0 = 16;
defparam sdpb_inst_182.BIT_WIDTH_1 = 16;
defparam sdpb_inst_182.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_182.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_182.RESET_MODE = "SYNC";

SDPB sdpb_inst_183 (
    .DO({sdpb_inst_183_dout_w[15:0],sdpb_inst_183_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_55}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_183}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_183.READ_MODE = 1'b0;
defparam sdpb_inst_183.BIT_WIDTH_0 = 16;
defparam sdpb_inst_183.BIT_WIDTH_1 = 16;
defparam sdpb_inst_183.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_183.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_183.RESET_MODE = "SYNC";

SDPB sdpb_inst_184 (
    .DO({sdpb_inst_184_dout_w[15:0],sdpb_inst_184_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_184}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_184.READ_MODE = 1'b0;
defparam sdpb_inst_184.BIT_WIDTH_0 = 16;
defparam sdpb_inst_184.BIT_WIDTH_1 = 16;
defparam sdpb_inst_184.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_184.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_184.RESET_MODE = "SYNC";

SDPB sdpb_inst_185 (
    .DO({sdpb_inst_185_dout_w[15:0],sdpb_inst_185_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_185}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_185.READ_MODE = 1'b0;
defparam sdpb_inst_185.BIT_WIDTH_0 = 16;
defparam sdpb_inst_185.BIT_WIDTH_1 = 16;
defparam sdpb_inst_185.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_185.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_185.RESET_MODE = "SYNC";

SDPB sdpb_inst_186 (
    .DO({sdpb_inst_186_dout_w[15:0],sdpb_inst_186_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_58}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_186}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_186.READ_MODE = 1'b0;
defparam sdpb_inst_186.BIT_WIDTH_0 = 16;
defparam sdpb_inst_186.BIT_WIDTH_1 = 16;
defparam sdpb_inst_186.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_186.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_186.RESET_MODE = "SYNC";

SDPB sdpb_inst_187 (
    .DO({sdpb_inst_187_dout_w[15:0],sdpb_inst_187_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_59}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_187}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_187.READ_MODE = 1'b0;
defparam sdpb_inst_187.BIT_WIDTH_0 = 16;
defparam sdpb_inst_187.BIT_WIDTH_1 = 16;
defparam sdpb_inst_187.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_187.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_187.RESET_MODE = "SYNC";

SDPB sdpb_inst_188 (
    .DO({sdpb_inst_188_dout_w[15:0],sdpb_inst_188_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_60}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_188}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_188.READ_MODE = 1'b0;
defparam sdpb_inst_188.BIT_WIDTH_0 = 16;
defparam sdpb_inst_188.BIT_WIDTH_1 = 16;
defparam sdpb_inst_188.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_188.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_188.RESET_MODE = "SYNC";

SDPB sdpb_inst_189 (
    .DO({sdpb_inst_189_dout_w[15:0],sdpb_inst_189_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_61}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_189}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_189.READ_MODE = 1'b0;
defparam sdpb_inst_189.BIT_WIDTH_0 = 16;
defparam sdpb_inst_189.BIT_WIDTH_1 = 16;
defparam sdpb_inst_189.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_189.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_189.RESET_MODE = "SYNC";

SDPB sdpb_inst_190 (
    .DO({sdpb_inst_190_dout_w[15:0],sdpb_inst_190_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_62}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_190}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_190.READ_MODE = 1'b0;
defparam sdpb_inst_190.BIT_WIDTH_0 = 16;
defparam sdpb_inst_190.BIT_WIDTH_1 = 16;
defparam sdpb_inst_190.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_190.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_190.RESET_MODE = "SYNC";

SDPB sdpb_inst_191 (
    .DO({sdpb_inst_191_dout_w[15:0],sdpb_inst_191_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_63}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_191}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_191.READ_MODE = 1'b0;
defparam sdpb_inst_191.BIT_WIDTH_0 = 16;
defparam sdpb_inst_191.BIT_WIDTH_1 = 16;
defparam sdpb_inst_191.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_191.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_191.RESET_MODE = "SYNC";

SDPB sdpb_inst_192 (
    .DO({sdpb_inst_192_dout_w[15:0],sdpb_inst_192_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_64}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_192}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_192.READ_MODE = 1'b0;
defparam sdpb_inst_192.BIT_WIDTH_0 = 16;
defparam sdpb_inst_192.BIT_WIDTH_1 = 16;
defparam sdpb_inst_192.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_192.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_192.RESET_MODE = "SYNC";

SDPB sdpb_inst_193 (
    .DO({sdpb_inst_193_dout_w[15:0],sdpb_inst_193_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_65}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_193}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_193.READ_MODE = 1'b0;
defparam sdpb_inst_193.BIT_WIDTH_0 = 16;
defparam sdpb_inst_193.BIT_WIDTH_1 = 16;
defparam sdpb_inst_193.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_193.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_193.RESET_MODE = "SYNC";

SDPB sdpb_inst_194 (
    .DO({sdpb_inst_194_dout_w[15:0],sdpb_inst_194_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_66}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_194}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_194.READ_MODE = 1'b0;
defparam sdpb_inst_194.BIT_WIDTH_0 = 16;
defparam sdpb_inst_194.BIT_WIDTH_1 = 16;
defparam sdpb_inst_194.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_194.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_194.RESET_MODE = "SYNC";

SDPB sdpb_inst_195 (
    .DO({sdpb_inst_195_dout_w[15:0],sdpb_inst_195_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_67}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_195}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_195.READ_MODE = 1'b0;
defparam sdpb_inst_195.BIT_WIDTH_0 = 16;
defparam sdpb_inst_195.BIT_WIDTH_1 = 16;
defparam sdpb_inst_195.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_195.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_195.RESET_MODE = "SYNC";

SDPB sdpb_inst_196 (
    .DO({sdpb_inst_196_dout_w[15:0],sdpb_inst_196_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_68}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_196}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_196.READ_MODE = 1'b0;
defparam sdpb_inst_196.BIT_WIDTH_0 = 16;
defparam sdpb_inst_196.BIT_WIDTH_1 = 16;
defparam sdpb_inst_196.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_196.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_196.RESET_MODE = "SYNC";

SDPB sdpb_inst_197 (
    .DO({sdpb_inst_197_dout_w[15:0],sdpb_inst_197_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_69}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_197}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_197.READ_MODE = 1'b0;
defparam sdpb_inst_197.BIT_WIDTH_0 = 16;
defparam sdpb_inst_197.BIT_WIDTH_1 = 16;
defparam sdpb_inst_197.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_197.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_197.RESET_MODE = "SYNC";

SDPB sdpb_inst_198 (
    .DO({sdpb_inst_198_dout_w[15:0],sdpb_inst_198_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_70}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_198}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_198.READ_MODE = 1'b0;
defparam sdpb_inst_198.BIT_WIDTH_0 = 16;
defparam sdpb_inst_198.BIT_WIDTH_1 = 16;
defparam sdpb_inst_198.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_198.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_198.RESET_MODE = "SYNC";

SDPB sdpb_inst_199 (
    .DO({sdpb_inst_199_dout_w[15:0],sdpb_inst_199_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_71}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_199}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_199.READ_MODE = 1'b0;
defparam sdpb_inst_199.BIT_WIDTH_0 = 16;
defparam sdpb_inst_199.BIT_WIDTH_1 = 16;
defparam sdpb_inst_199.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_199.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_199.RESET_MODE = "SYNC";

SDPB sdpb_inst_200 (
    .DO({sdpb_inst_200_dout_w[15:0],sdpb_inst_200_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_72}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_200}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_200.READ_MODE = 1'b0;
defparam sdpb_inst_200.BIT_WIDTH_0 = 16;
defparam sdpb_inst_200.BIT_WIDTH_1 = 16;
defparam sdpb_inst_200.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_200.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_200.RESET_MODE = "SYNC";

SDPB sdpb_inst_201 (
    .DO({sdpb_inst_201_dout_w[15:0],sdpb_inst_201_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_73}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_201}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_201.READ_MODE = 1'b0;
defparam sdpb_inst_201.BIT_WIDTH_0 = 16;
defparam sdpb_inst_201.BIT_WIDTH_1 = 16;
defparam sdpb_inst_201.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_201.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_201.RESET_MODE = "SYNC";

SDPB sdpb_inst_202 (
    .DO({sdpb_inst_202_dout_w[15:0],sdpb_inst_202_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_74}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_202}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_202.READ_MODE = 1'b0;
defparam sdpb_inst_202.BIT_WIDTH_0 = 16;
defparam sdpb_inst_202.BIT_WIDTH_1 = 16;
defparam sdpb_inst_202.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_202.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_202.RESET_MODE = "SYNC";

SDPB sdpb_inst_203 (
    .DO({sdpb_inst_203_dout_w[15:0],sdpb_inst_203_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_75}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_203}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_203.READ_MODE = 1'b0;
defparam sdpb_inst_203.BIT_WIDTH_0 = 16;
defparam sdpb_inst_203.BIT_WIDTH_1 = 16;
defparam sdpb_inst_203.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_203.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_203.RESET_MODE = "SYNC";

SDPB sdpb_inst_204 (
    .DO({sdpb_inst_204_dout_w[15:0],sdpb_inst_204_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_76}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_204}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_204.READ_MODE = 1'b0;
defparam sdpb_inst_204.BIT_WIDTH_0 = 16;
defparam sdpb_inst_204.BIT_WIDTH_1 = 16;
defparam sdpb_inst_204.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_204.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_204.RESET_MODE = "SYNC";

SDPB sdpb_inst_205 (
    .DO({sdpb_inst_205_dout_w[15:0],sdpb_inst_205_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_77}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_205}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_205.READ_MODE = 1'b0;
defparam sdpb_inst_205.BIT_WIDTH_0 = 16;
defparam sdpb_inst_205.BIT_WIDTH_1 = 16;
defparam sdpb_inst_205.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_205.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_205.RESET_MODE = "SYNC";

SDPB sdpb_inst_206 (
    .DO({sdpb_inst_206_dout_w[15:0],sdpb_inst_206_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_78}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_206}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_206.READ_MODE = 1'b0;
defparam sdpb_inst_206.BIT_WIDTH_0 = 16;
defparam sdpb_inst_206.BIT_WIDTH_1 = 16;
defparam sdpb_inst_206.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_206.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_206.RESET_MODE = "SYNC";

SDPB sdpb_inst_207 (
    .DO({sdpb_inst_207_dout_w[15:0],sdpb_inst_207_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_79}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_207}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_207.READ_MODE = 1'b0;
defparam sdpb_inst_207.BIT_WIDTH_0 = 16;
defparam sdpb_inst_207.BIT_WIDTH_1 = 16;
defparam sdpb_inst_207.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_207.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_207.RESET_MODE = "SYNC";

SDPB sdpb_inst_208 (
    .DO({sdpb_inst_208_dout_w[15:0],sdpb_inst_208_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_80}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_208}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_208.READ_MODE = 1'b0;
defparam sdpb_inst_208.BIT_WIDTH_0 = 16;
defparam sdpb_inst_208.BIT_WIDTH_1 = 16;
defparam sdpb_inst_208.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_208.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_208.RESET_MODE = "SYNC";

SDPB sdpb_inst_209 (
    .DO({sdpb_inst_209_dout_w[15:0],sdpb_inst_209_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_81}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_209}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_209.READ_MODE = 1'b0;
defparam sdpb_inst_209.BIT_WIDTH_0 = 16;
defparam sdpb_inst_209.BIT_WIDTH_1 = 16;
defparam sdpb_inst_209.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_209.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_209.RESET_MODE = "SYNC";

SDPB sdpb_inst_210 (
    .DO({sdpb_inst_210_dout_w[15:0],sdpb_inst_210_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_82}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_210}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_210.READ_MODE = 1'b0;
defparam sdpb_inst_210.BIT_WIDTH_0 = 16;
defparam sdpb_inst_210.BIT_WIDTH_1 = 16;
defparam sdpb_inst_210.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_210.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_210.RESET_MODE = "SYNC";

SDPB sdpb_inst_211 (
    .DO({sdpb_inst_211_dout_w[15:0],sdpb_inst_211_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_83}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_211}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_211.READ_MODE = 1'b0;
defparam sdpb_inst_211.BIT_WIDTH_0 = 16;
defparam sdpb_inst_211.BIT_WIDTH_1 = 16;
defparam sdpb_inst_211.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_211.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_211.RESET_MODE = "SYNC";

SDPB sdpb_inst_212 (
    .DO({sdpb_inst_212_dout_w[15:0],sdpb_inst_212_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_84}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_212}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_212.READ_MODE = 1'b0;
defparam sdpb_inst_212.BIT_WIDTH_0 = 16;
defparam sdpb_inst_212.BIT_WIDTH_1 = 16;
defparam sdpb_inst_212.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_212.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_212.RESET_MODE = "SYNC";

SDPB sdpb_inst_213 (
    .DO({sdpb_inst_213_dout_w[15:0],sdpb_inst_213_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_85}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_213}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_213.READ_MODE = 1'b0;
defparam sdpb_inst_213.BIT_WIDTH_0 = 16;
defparam sdpb_inst_213.BIT_WIDTH_1 = 16;
defparam sdpb_inst_213.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_213.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_213.RESET_MODE = "SYNC";

SDPB sdpb_inst_214 (
    .DO({sdpb_inst_214_dout_w[15:0],sdpb_inst_214_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_86}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_214}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_214.READ_MODE = 1'b0;
defparam sdpb_inst_214.BIT_WIDTH_0 = 16;
defparam sdpb_inst_214.BIT_WIDTH_1 = 16;
defparam sdpb_inst_214.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_214.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_214.RESET_MODE = "SYNC";

SDPB sdpb_inst_215 (
    .DO({sdpb_inst_215_dout_w[15:0],sdpb_inst_215_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_87}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_215}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_215.READ_MODE = 1'b0;
defparam sdpb_inst_215.BIT_WIDTH_0 = 16;
defparam sdpb_inst_215.BIT_WIDTH_1 = 16;
defparam sdpb_inst_215.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_215.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_215.RESET_MODE = "SYNC";

SDPB sdpb_inst_216 (
    .DO({sdpb_inst_216_dout_w[15:0],sdpb_inst_216_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_88}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_216}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_216.READ_MODE = 1'b0;
defparam sdpb_inst_216.BIT_WIDTH_0 = 16;
defparam sdpb_inst_216.BIT_WIDTH_1 = 16;
defparam sdpb_inst_216.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_216.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_216.RESET_MODE = "SYNC";

SDPB sdpb_inst_217 (
    .DO({sdpb_inst_217_dout_w[15:0],sdpb_inst_217_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_89}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_217}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_217.READ_MODE = 1'b0;
defparam sdpb_inst_217.BIT_WIDTH_0 = 16;
defparam sdpb_inst_217.BIT_WIDTH_1 = 16;
defparam sdpb_inst_217.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_217.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_217.RESET_MODE = "SYNC";

SDPB sdpb_inst_218 (
    .DO({sdpb_inst_218_dout_w[15:0],sdpb_inst_218_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_90}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_218}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_218.READ_MODE = 1'b0;
defparam sdpb_inst_218.BIT_WIDTH_0 = 16;
defparam sdpb_inst_218.BIT_WIDTH_1 = 16;
defparam sdpb_inst_218.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_218.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_218.RESET_MODE = "SYNC";

SDPB sdpb_inst_219 (
    .DO({sdpb_inst_219_dout_w[15:0],sdpb_inst_219_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_91}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_219}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_219.READ_MODE = 1'b0;
defparam sdpb_inst_219.BIT_WIDTH_0 = 16;
defparam sdpb_inst_219.BIT_WIDTH_1 = 16;
defparam sdpb_inst_219.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_219.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_219.RESET_MODE = "SYNC";

SDPB sdpb_inst_220 (
    .DO({sdpb_inst_220_dout_w[15:0],sdpb_inst_220_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_92}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_220}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_220.READ_MODE = 1'b0;
defparam sdpb_inst_220.BIT_WIDTH_0 = 16;
defparam sdpb_inst_220.BIT_WIDTH_1 = 16;
defparam sdpb_inst_220.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_220.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_220.RESET_MODE = "SYNC";

SDPB sdpb_inst_221 (
    .DO({sdpb_inst_221_dout_w[15:0],sdpb_inst_221_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_93}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_221}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_221.READ_MODE = 1'b0;
defparam sdpb_inst_221.BIT_WIDTH_0 = 16;
defparam sdpb_inst_221.BIT_WIDTH_1 = 16;
defparam sdpb_inst_221.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_221.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_221.RESET_MODE = "SYNC";

SDPB sdpb_inst_222 (
    .DO({sdpb_inst_222_dout_w[15:0],sdpb_inst_222_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_94}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_222}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_222.READ_MODE = 1'b0;
defparam sdpb_inst_222.BIT_WIDTH_0 = 16;
defparam sdpb_inst_222.BIT_WIDTH_1 = 16;
defparam sdpb_inst_222.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_222.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_222.RESET_MODE = "SYNC";

SDPB sdpb_inst_223 (
    .DO({sdpb_inst_223_dout_w[15:0],sdpb_inst_223_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_95}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_223}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_223.READ_MODE = 1'b0;
defparam sdpb_inst_223.BIT_WIDTH_0 = 16;
defparam sdpb_inst_223.BIT_WIDTH_1 = 16;
defparam sdpb_inst_223.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_223.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_223.RESET_MODE = "SYNC";

SDPB sdpb_inst_224 (
    .DO({sdpb_inst_224_dout_w[15:0],sdpb_inst_224_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_96}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_224}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_224.READ_MODE = 1'b0;
defparam sdpb_inst_224.BIT_WIDTH_0 = 16;
defparam sdpb_inst_224.BIT_WIDTH_1 = 16;
defparam sdpb_inst_224.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_224.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_224.RESET_MODE = "SYNC";

SDPB sdpb_inst_225 (
    .DO({sdpb_inst_225_dout_w[15:0],sdpb_inst_225_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_97}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_225}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_225.READ_MODE = 1'b0;
defparam sdpb_inst_225.BIT_WIDTH_0 = 16;
defparam sdpb_inst_225.BIT_WIDTH_1 = 16;
defparam sdpb_inst_225.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_225.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_225.RESET_MODE = "SYNC";

SDPB sdpb_inst_226 (
    .DO({sdpb_inst_226_dout_w[15:0],sdpb_inst_226_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_98}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_226}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_226.READ_MODE = 1'b0;
defparam sdpb_inst_226.BIT_WIDTH_0 = 16;
defparam sdpb_inst_226.BIT_WIDTH_1 = 16;
defparam sdpb_inst_226.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_226.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_226.RESET_MODE = "SYNC";

SDPB sdpb_inst_227 (
    .DO({sdpb_inst_227_dout_w[15:0],sdpb_inst_227_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_99}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_227}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_227.READ_MODE = 1'b0;
defparam sdpb_inst_227.BIT_WIDTH_0 = 16;
defparam sdpb_inst_227.BIT_WIDTH_1 = 16;
defparam sdpb_inst_227.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_227.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_227.RESET_MODE = "SYNC";

SDPB sdpb_inst_228 (
    .DO({sdpb_inst_228_dout_w[15:0],sdpb_inst_228_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_100}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_228}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_228.READ_MODE = 1'b0;
defparam sdpb_inst_228.BIT_WIDTH_0 = 16;
defparam sdpb_inst_228.BIT_WIDTH_1 = 16;
defparam sdpb_inst_228.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_228.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_228.RESET_MODE = "SYNC";

SDPB sdpb_inst_229 (
    .DO({sdpb_inst_229_dout_w[15:0],sdpb_inst_229_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_101}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_229}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_229.READ_MODE = 1'b0;
defparam sdpb_inst_229.BIT_WIDTH_0 = 16;
defparam sdpb_inst_229.BIT_WIDTH_1 = 16;
defparam sdpb_inst_229.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_229.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_229.RESET_MODE = "SYNC";

SDPB sdpb_inst_230 (
    .DO({sdpb_inst_230_dout_w[15:0],sdpb_inst_230_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_102}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_230}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_230.READ_MODE = 1'b0;
defparam sdpb_inst_230.BIT_WIDTH_0 = 16;
defparam sdpb_inst_230.BIT_WIDTH_1 = 16;
defparam sdpb_inst_230.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_230.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_230.RESET_MODE = "SYNC";

SDPB sdpb_inst_231 (
    .DO({sdpb_inst_231_dout_w[15:0],sdpb_inst_231_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_103}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_231}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_231.READ_MODE = 1'b0;
defparam sdpb_inst_231.BIT_WIDTH_0 = 16;
defparam sdpb_inst_231.BIT_WIDTH_1 = 16;
defparam sdpb_inst_231.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_231.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_231.RESET_MODE = "SYNC";

SDPB sdpb_inst_232 (
    .DO({sdpb_inst_232_dout_w[15:0],sdpb_inst_232_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_104}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_232}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_232.READ_MODE = 1'b0;
defparam sdpb_inst_232.BIT_WIDTH_0 = 16;
defparam sdpb_inst_232.BIT_WIDTH_1 = 16;
defparam sdpb_inst_232.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_232.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_232.RESET_MODE = "SYNC";

SDPB sdpb_inst_233 (
    .DO({sdpb_inst_233_dout_w[15:0],sdpb_inst_233_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_105}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_233}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_233.READ_MODE = 1'b0;
defparam sdpb_inst_233.BIT_WIDTH_0 = 16;
defparam sdpb_inst_233.BIT_WIDTH_1 = 16;
defparam sdpb_inst_233.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_233.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_233.RESET_MODE = "SYNC";

SDPB sdpb_inst_234 (
    .DO({sdpb_inst_234_dout_w[15:0],sdpb_inst_234_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_106}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_234}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_234.READ_MODE = 1'b0;
defparam sdpb_inst_234.BIT_WIDTH_0 = 16;
defparam sdpb_inst_234.BIT_WIDTH_1 = 16;
defparam sdpb_inst_234.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_234.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_234.RESET_MODE = "SYNC";

SDPB sdpb_inst_235 (
    .DO({sdpb_inst_235_dout_w[15:0],sdpb_inst_235_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_107}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_235}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_235.READ_MODE = 1'b0;
defparam sdpb_inst_235.BIT_WIDTH_0 = 16;
defparam sdpb_inst_235.BIT_WIDTH_1 = 16;
defparam sdpb_inst_235.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_235.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_235.RESET_MODE = "SYNC";

SDPB sdpb_inst_236 (
    .DO({sdpb_inst_236_dout_w[15:0],sdpb_inst_236_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_108}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_236}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_236.READ_MODE = 1'b0;
defparam sdpb_inst_236.BIT_WIDTH_0 = 16;
defparam sdpb_inst_236.BIT_WIDTH_1 = 16;
defparam sdpb_inst_236.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_236.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_236.RESET_MODE = "SYNC";

SDPB sdpb_inst_237 (
    .DO({sdpb_inst_237_dout_w[15:0],sdpb_inst_237_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_109}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_237}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_237.READ_MODE = 1'b0;
defparam sdpb_inst_237.BIT_WIDTH_0 = 16;
defparam sdpb_inst_237.BIT_WIDTH_1 = 16;
defparam sdpb_inst_237.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_237.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_237.RESET_MODE = "SYNC";

SDPB sdpb_inst_238 (
    .DO({sdpb_inst_238_dout_w[15:0],sdpb_inst_238_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_110}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_238}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_238.READ_MODE = 1'b0;
defparam sdpb_inst_238.BIT_WIDTH_0 = 16;
defparam sdpb_inst_238.BIT_WIDTH_1 = 16;
defparam sdpb_inst_238.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_238.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_238.RESET_MODE = "SYNC";

SDPB sdpb_inst_239 (
    .DO({sdpb_inst_239_dout_w[15:0],sdpb_inst_239_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_111}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_239}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_239.READ_MODE = 1'b0;
defparam sdpb_inst_239.BIT_WIDTH_0 = 16;
defparam sdpb_inst_239.BIT_WIDTH_1 = 16;
defparam sdpb_inst_239.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_239.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_239.RESET_MODE = "SYNC";

SDPB sdpb_inst_240 (
    .DO({sdpb_inst_240_dout_w[15:0],sdpb_inst_240_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_112}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_240}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_240.READ_MODE = 1'b0;
defparam sdpb_inst_240.BIT_WIDTH_0 = 16;
defparam sdpb_inst_240.BIT_WIDTH_1 = 16;
defparam sdpb_inst_240.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_240.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_240.RESET_MODE = "SYNC";

SDPB sdpb_inst_241 (
    .DO({sdpb_inst_241_dout_w[15:0],sdpb_inst_241_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_113}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_241}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_241.READ_MODE = 1'b0;
defparam sdpb_inst_241.BIT_WIDTH_0 = 16;
defparam sdpb_inst_241.BIT_WIDTH_1 = 16;
defparam sdpb_inst_241.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_241.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_241.RESET_MODE = "SYNC";

SDPB sdpb_inst_242 (
    .DO({sdpb_inst_242_dout_w[15:0],sdpb_inst_242_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_114}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_242}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_242.READ_MODE = 1'b0;
defparam sdpb_inst_242.BIT_WIDTH_0 = 16;
defparam sdpb_inst_242.BIT_WIDTH_1 = 16;
defparam sdpb_inst_242.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_242.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_242.RESET_MODE = "SYNC";

SDPB sdpb_inst_243 (
    .DO({sdpb_inst_243_dout_w[15:0],sdpb_inst_243_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_115}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_243}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_243.READ_MODE = 1'b0;
defparam sdpb_inst_243.BIT_WIDTH_0 = 16;
defparam sdpb_inst_243.BIT_WIDTH_1 = 16;
defparam sdpb_inst_243.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_243.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_243.RESET_MODE = "SYNC";

SDPB sdpb_inst_244 (
    .DO({sdpb_inst_244_dout_w[15:0],sdpb_inst_244_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_116}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_244}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_244.READ_MODE = 1'b0;
defparam sdpb_inst_244.BIT_WIDTH_0 = 16;
defparam sdpb_inst_244.BIT_WIDTH_1 = 16;
defparam sdpb_inst_244.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_244.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_244.RESET_MODE = "SYNC";

SDPB sdpb_inst_245 (
    .DO({sdpb_inst_245_dout_w[15:0],sdpb_inst_245_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_117}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_245}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_245.READ_MODE = 1'b0;
defparam sdpb_inst_245.BIT_WIDTH_0 = 16;
defparam sdpb_inst_245.BIT_WIDTH_1 = 16;
defparam sdpb_inst_245.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_245.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_245.RESET_MODE = "SYNC";

SDPB sdpb_inst_246 (
    .DO({sdpb_inst_246_dout_w[15:0],sdpb_inst_246_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_118}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_246}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_246.READ_MODE = 1'b0;
defparam sdpb_inst_246.BIT_WIDTH_0 = 16;
defparam sdpb_inst_246.BIT_WIDTH_1 = 16;
defparam sdpb_inst_246.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_246.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_246.RESET_MODE = "SYNC";

SDPB sdpb_inst_247 (
    .DO({sdpb_inst_247_dout_w[15:0],sdpb_inst_247_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_119}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_247}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_247.READ_MODE = 1'b0;
defparam sdpb_inst_247.BIT_WIDTH_0 = 16;
defparam sdpb_inst_247.BIT_WIDTH_1 = 16;
defparam sdpb_inst_247.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_247.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_247.RESET_MODE = "SYNC";

SDPB sdpb_inst_248 (
    .DO({sdpb_inst_248_dout_w[15:0],sdpb_inst_248_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_120}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_248}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_248.READ_MODE = 1'b0;
defparam sdpb_inst_248.BIT_WIDTH_0 = 16;
defparam sdpb_inst_248.BIT_WIDTH_1 = 16;
defparam sdpb_inst_248.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_248.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_248.RESET_MODE = "SYNC";

SDPB sdpb_inst_249 (
    .DO({sdpb_inst_249_dout_w[15:0],sdpb_inst_249_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_121}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_249}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_249.READ_MODE = 1'b0;
defparam sdpb_inst_249.BIT_WIDTH_0 = 16;
defparam sdpb_inst_249.BIT_WIDTH_1 = 16;
defparam sdpb_inst_249.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_249.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_249.RESET_MODE = "SYNC";

SDPB sdpb_inst_250 (
    .DO({sdpb_inst_250_dout_w[15:0],sdpb_inst_250_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_122}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_250}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_250.READ_MODE = 1'b0;
defparam sdpb_inst_250.BIT_WIDTH_0 = 16;
defparam sdpb_inst_250.BIT_WIDTH_1 = 16;
defparam sdpb_inst_250.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_250.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_250.RESET_MODE = "SYNC";

SDPB sdpb_inst_251 (
    .DO({sdpb_inst_251_dout_w[15:0],sdpb_inst_251_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_123}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_251}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_251.READ_MODE = 1'b0;
defparam sdpb_inst_251.BIT_WIDTH_0 = 16;
defparam sdpb_inst_251.BIT_WIDTH_1 = 16;
defparam sdpb_inst_251.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_251.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_251.RESET_MODE = "SYNC";

SDPB sdpb_inst_252 (
    .DO({sdpb_inst_252_dout_w[15:0],sdpb_inst_252_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_124}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_252}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_252.READ_MODE = 1'b0;
defparam sdpb_inst_252.BIT_WIDTH_0 = 16;
defparam sdpb_inst_252.BIT_WIDTH_1 = 16;
defparam sdpb_inst_252.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_252.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_252.RESET_MODE = "SYNC";

SDPB sdpb_inst_253 (
    .DO({sdpb_inst_253_dout_w[15:0],sdpb_inst_253_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_125}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_253}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_253.READ_MODE = 1'b0;
defparam sdpb_inst_253.BIT_WIDTH_0 = 16;
defparam sdpb_inst_253.BIT_WIDTH_1 = 16;
defparam sdpb_inst_253.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_253.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_253.RESET_MODE = "SYNC";

SDPB sdpb_inst_254 (
    .DO({sdpb_inst_254_dout_w[15:0],sdpb_inst_254_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_126}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_254}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_254.READ_MODE = 1'b0;
defparam sdpb_inst_254.BIT_WIDTH_0 = 16;
defparam sdpb_inst_254.BIT_WIDTH_1 = 16;
defparam sdpb_inst_254.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_254.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_254.RESET_MODE = "SYNC";

SDPB sdpb_inst_255 (
    .DO({sdpb_inst_255_dout_w[15:0],sdpb_inst_255_dout[31:16]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_127}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_255}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_255.READ_MODE = 1'b0;
defparam sdpb_inst_255.BIT_WIDTH_0 = 16;
defparam sdpb_inst_255.BIT_WIDTH_1 = 16;
defparam sdpb_inst_255.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_255.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_255.RESET_MODE = "SYNC";

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[16]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_6 (
  .Q(dff_q_6),
  .D(adb[10]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sdpb_inst_2_dout[0]),
  .I1(sdpb_inst_3_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sdpb_inst_4_dout[0]),
  .I1(sdpb_inst_5_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sdpb_inst_6_dout[0]),
  .I1(sdpb_inst_7_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sdpb_inst_8_dout[0]),
  .I1(sdpb_inst_9_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sdpb_inst_10_dout[0]),
  .I1(sdpb_inst_11_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sdpb_inst_12_dout[0]),
  .I1(sdpb_inst_13_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(sdpb_inst_14_dout[0]),
  .I1(sdpb_inst_15_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sdpb_inst_16_dout[0]),
  .I1(sdpb_inst_17_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(sdpb_inst_18_dout[0]),
  .I1(sdpb_inst_19_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(sdpb_inst_20_dout[0]),
  .I1(sdpb_inst_21_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(sdpb_inst_22_dout[0]),
  .I1(sdpb_inst_23_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(sdpb_inst_24_dout[0]),
  .I1(sdpb_inst_25_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(sdpb_inst_26_dout[0]),
  .I1(sdpb_inst_27_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(sdpb_inst_28_dout[0]),
  .I1(sdpb_inst_29_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sdpb_inst_30_dout[0]),
  .I1(sdpb_inst_31_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sdpb_inst_32_dout[0]),
  .I1(sdpb_inst_33_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(sdpb_inst_34_dout[0]),
  .I1(sdpb_inst_35_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(sdpb_inst_36_dout[0]),
  .I1(sdpb_inst_37_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(sdpb_inst_38_dout[0]),
  .I1(sdpb_inst_39_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(sdpb_inst_40_dout[0]),
  .I1(sdpb_inst_41_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sdpb_inst_42_dout[0]),
  .I1(sdpb_inst_43_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(sdpb_inst_44_dout[0]),
  .I1(sdpb_inst_45_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(sdpb_inst_46_dout[0]),
  .I1(sdpb_inst_47_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(sdpb_inst_48_dout[0]),
  .I1(sdpb_inst_49_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(sdpb_inst_50_dout[0]),
  .I1(sdpb_inst_51_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(sdpb_inst_52_dout[0]),
  .I1(sdpb_inst_53_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(sdpb_inst_54_dout[0]),
  .I1(sdpb_inst_55_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(sdpb_inst_56_dout[0]),
  .I1(sdpb_inst_57_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(sdpb_inst_58_dout[0]),
  .I1(sdpb_inst_59_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(sdpb_inst_60_dout[0]),
  .I1(sdpb_inst_61_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(sdpb_inst_62_dout[0]),
  .I1(sdpb_inst_63_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(sdpb_inst_64_dout[0]),
  .I1(sdpb_inst_65_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sdpb_inst_66_dout[0]),
  .I1(sdpb_inst_67_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(sdpb_inst_68_dout[0]),
  .I1(sdpb_inst_69_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(sdpb_inst_70_dout[0]),
  .I1(sdpb_inst_71_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sdpb_inst_72_dout[0]),
  .I1(sdpb_inst_73_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(sdpb_inst_74_dout[0]),
  .I1(sdpb_inst_75_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(sdpb_inst_76_dout[0]),
  .I1(sdpb_inst_77_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(sdpb_inst_78_dout[0]),
  .I1(sdpb_inst_79_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(sdpb_inst_80_dout[0]),
  .I1(sdpb_inst_81_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(sdpb_inst_82_dout[0]),
  .I1(sdpb_inst_83_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(sdpb_inst_84_dout[0]),
  .I1(sdpb_inst_85_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(sdpb_inst_86_dout[0]),
  .I1(sdpb_inst_87_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(sdpb_inst_88_dout[0]),
  .I1(sdpb_inst_89_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sdpb_inst_90_dout[0]),
  .I1(sdpb_inst_91_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sdpb_inst_92_dout[0]),
  .I1(sdpb_inst_93_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(sdpb_inst_94_dout[0]),
  .I1(sdpb_inst_95_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(sdpb_inst_96_dout[0]),
  .I1(sdpb_inst_97_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(sdpb_inst_98_dout[0]),
  .I1(sdpb_inst_99_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(sdpb_inst_100_dout[0]),
  .I1(sdpb_inst_101_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(sdpb_inst_102_dout[0]),
  .I1(sdpb_inst_103_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(sdpb_inst_104_dout[0]),
  .I1(sdpb_inst_105_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(sdpb_inst_106_dout[0]),
  .I1(sdpb_inst_107_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(sdpb_inst_108_dout[0]),
  .I1(sdpb_inst_109_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(sdpb_inst_110_dout[0]),
  .I1(sdpb_inst_111_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(sdpb_inst_112_dout[0]),
  .I1(sdpb_inst_113_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(sdpb_inst_114_dout[0]),
  .I1(sdpb_inst_115_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(sdpb_inst_116_dout[0]),
  .I1(sdpb_inst_117_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(sdpb_inst_118_dout[0]),
  .I1(sdpb_inst_119_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(sdpb_inst_120_dout[0]),
  .I1(sdpb_inst_121_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(sdpb_inst_122_dout[0]),
  .I1(sdpb_inst_123_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(sdpb_inst_124_dout[0]),
  .I1(sdpb_inst_125_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sdpb_inst_126_dout[0]),
  .I1(sdpb_inst_127_dout[0]),
  .S0(dff_q_6)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_5)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_5)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_5)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_5)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_5)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_5)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_5)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_5)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_5)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_5)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(dff_q_5)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(dff_q_5)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(dff_q_5)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(dff_q_5)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_5)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_5)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_5)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(dff_q_5)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(dff_q_5)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_5)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_5)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_5)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(dff_q_5)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(dff_q_5)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_48),
  .I1(mux_o_49),
  .S0(dff_q_5)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_50),
  .I1(mux_o_51),
  .S0(dff_q_5)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_52),
  .I1(mux_o_53),
  .S0(dff_q_5)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(dff_q_5)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(dff_q_5)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(dff_q_5)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_5)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_5)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(dff_q_4)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_4)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(dff_q_4)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_4)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_4)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(dff_q_4)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_76),
  .I1(mux_o_77),
  .S0(dff_q_4)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_78),
  .I1(mux_o_79),
  .S0(dff_q_4)
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(mux_o_80),
  .I1(mux_o_81),
  .S0(dff_q_4)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(mux_o_82),
  .I1(mux_o_83),
  .S0(dff_q_4)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(dff_q_4)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_4)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_4)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_4)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_4)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_4)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_3)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_3)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_3)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_104),
  .I1(mux_o_105),
  .S0(dff_q_3)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_106),
  .I1(mux_o_107),
  .S0(dff_q_3)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(dff_q_3)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_110),
  .I1(mux_o_111),
  .S0(dff_q_3)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(dff_q_2)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(dff_q_2)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_118),
  .I1(mux_o_119),
  .S0(dff_q_2)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(dff_q_1)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(dff_q_1)
);
MUX2 mux_inst_126 (
  .O(dout[0]),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(dff_q_0)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(sdpb_inst_0_dout[1]),
  .I1(sdpb_inst_1_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(sdpb_inst_2_dout[1]),
  .I1(sdpb_inst_3_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(sdpb_inst_4_dout[1]),
  .I1(sdpb_inst_5_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(sdpb_inst_6_dout[1]),
  .I1(sdpb_inst_7_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(sdpb_inst_8_dout[1]),
  .I1(sdpb_inst_9_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(sdpb_inst_10_dout[1]),
  .I1(sdpb_inst_11_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(sdpb_inst_12_dout[1]),
  .I1(sdpb_inst_13_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(sdpb_inst_14_dout[1]),
  .I1(sdpb_inst_15_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(sdpb_inst_16_dout[1]),
  .I1(sdpb_inst_17_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sdpb_inst_18_dout[1]),
  .I1(sdpb_inst_19_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(sdpb_inst_20_dout[1]),
  .I1(sdpb_inst_21_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(sdpb_inst_22_dout[1]),
  .I1(sdpb_inst_23_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(sdpb_inst_24_dout[1]),
  .I1(sdpb_inst_25_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(sdpb_inst_26_dout[1]),
  .I1(sdpb_inst_27_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(sdpb_inst_28_dout[1]),
  .I1(sdpb_inst_29_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(sdpb_inst_30_dout[1]),
  .I1(sdpb_inst_31_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(sdpb_inst_32_dout[1]),
  .I1(sdpb_inst_33_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(sdpb_inst_34_dout[1]),
  .I1(sdpb_inst_35_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(sdpb_inst_36_dout[1]),
  .I1(sdpb_inst_37_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(sdpb_inst_38_dout[1]),
  .I1(sdpb_inst_39_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(sdpb_inst_40_dout[1]),
  .I1(sdpb_inst_41_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(sdpb_inst_42_dout[1]),
  .I1(sdpb_inst_43_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(sdpb_inst_44_dout[1]),
  .I1(sdpb_inst_45_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(sdpb_inst_46_dout[1]),
  .I1(sdpb_inst_47_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(sdpb_inst_48_dout[1]),
  .I1(sdpb_inst_49_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(sdpb_inst_50_dout[1]),
  .I1(sdpb_inst_51_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(sdpb_inst_52_dout[1]),
  .I1(sdpb_inst_53_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(sdpb_inst_54_dout[1]),
  .I1(sdpb_inst_55_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(sdpb_inst_56_dout[1]),
  .I1(sdpb_inst_57_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(sdpb_inst_58_dout[1]),
  .I1(sdpb_inst_59_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(sdpb_inst_60_dout[1]),
  .I1(sdpb_inst_61_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(sdpb_inst_62_dout[1]),
  .I1(sdpb_inst_63_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(sdpb_inst_64_dout[1]),
  .I1(sdpb_inst_65_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(sdpb_inst_66_dout[1]),
  .I1(sdpb_inst_67_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(sdpb_inst_68_dout[1]),
  .I1(sdpb_inst_69_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(sdpb_inst_70_dout[1]),
  .I1(sdpb_inst_71_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(sdpb_inst_72_dout[1]),
  .I1(sdpb_inst_73_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(sdpb_inst_74_dout[1]),
  .I1(sdpb_inst_75_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(sdpb_inst_76_dout[1]),
  .I1(sdpb_inst_77_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(sdpb_inst_78_dout[1]),
  .I1(sdpb_inst_79_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(sdpb_inst_80_dout[1]),
  .I1(sdpb_inst_81_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(sdpb_inst_82_dout[1]),
  .I1(sdpb_inst_83_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(sdpb_inst_84_dout[1]),
  .I1(sdpb_inst_85_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(sdpb_inst_86_dout[1]),
  .I1(sdpb_inst_87_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(sdpb_inst_88_dout[1]),
  .I1(sdpb_inst_89_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(sdpb_inst_90_dout[1]),
  .I1(sdpb_inst_91_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(sdpb_inst_92_dout[1]),
  .I1(sdpb_inst_93_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(sdpb_inst_94_dout[1]),
  .I1(sdpb_inst_95_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(sdpb_inst_96_dout[1]),
  .I1(sdpb_inst_97_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(sdpb_inst_98_dout[1]),
  .I1(sdpb_inst_99_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(sdpb_inst_100_dout[1]),
  .I1(sdpb_inst_101_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(sdpb_inst_102_dout[1]),
  .I1(sdpb_inst_103_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(sdpb_inst_104_dout[1]),
  .I1(sdpb_inst_105_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(sdpb_inst_106_dout[1]),
  .I1(sdpb_inst_107_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(sdpb_inst_108_dout[1]),
  .I1(sdpb_inst_109_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(sdpb_inst_110_dout[1]),
  .I1(sdpb_inst_111_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(sdpb_inst_112_dout[1]),
  .I1(sdpb_inst_113_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(sdpb_inst_114_dout[1]),
  .I1(sdpb_inst_115_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(sdpb_inst_116_dout[1]),
  .I1(sdpb_inst_117_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(sdpb_inst_118_dout[1]),
  .I1(sdpb_inst_119_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(sdpb_inst_120_dout[1]),
  .I1(sdpb_inst_121_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(sdpb_inst_122_dout[1]),
  .I1(sdpb_inst_123_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(sdpb_inst_124_dout[1]),
  .I1(sdpb_inst_125_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(sdpb_inst_126_dout[1]),
  .I1(sdpb_inst_127_dout[1]),
  .S0(dff_q_6)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_127),
  .I1(mux_o_128),
  .S0(dff_q_5)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_129),
  .I1(mux_o_130),
  .S0(dff_q_5)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(dff_q_5)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_5)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_5)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_5)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(dff_q_5)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(dff_q_5)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(mux_o_143),
  .I1(mux_o_144),
  .S0(dff_q_5)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(dff_q_5)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_5)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(dff_q_5)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_151),
  .I1(mux_o_152),
  .S0(dff_q_5)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_153),
  .I1(mux_o_154),
  .S0(dff_q_5)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_155),
  .I1(mux_o_156),
  .S0(dff_q_5)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_157),
  .I1(mux_o_158),
  .S0(dff_q_5)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_159),
  .I1(mux_o_160),
  .S0(dff_q_5)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_5)
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(dff_q_5)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_5)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(dff_q_5)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(dff_q_5)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_5)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_5)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_5)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_5)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_5)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_5)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_5)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_185),
  .I1(mux_o_186),
  .S0(dff_q_5)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_187),
  .I1(mux_o_188),
  .S0(dff_q_5)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_5)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(dff_q_4)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(dff_q_4)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(dff_q_4)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(dff_q_4)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(dff_q_4)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_4)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_4)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_4)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_4)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(mux_o_209),
  .I1(mux_o_210),
  .S0(dff_q_4)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_211),
  .I1(mux_o_212),
  .S0(dff_q_4)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_213),
  .I1(mux_o_214),
  .S0(dff_q_4)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_215),
  .I1(mux_o_216),
  .S0(dff_q_4)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_4)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_4)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_4)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(dff_q_3)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_3)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_3)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_3)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_3)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_3)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_2)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(dff_q_2)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(dff_q_2)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_2)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_247),
  .I1(mux_o_248),
  .S0(dff_q_1)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(dff_q_1)
);
MUX2 mux_inst_253 (
  .O(dout[1]),
  .I0(mux_o_251),
  .I1(mux_o_252),
  .S0(dff_q_0)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(sdpb_inst_0_dout[2]),
  .I1(sdpb_inst_1_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(sdpb_inst_2_dout[2]),
  .I1(sdpb_inst_3_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(sdpb_inst_4_dout[2]),
  .I1(sdpb_inst_5_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(sdpb_inst_6_dout[2]),
  .I1(sdpb_inst_7_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(sdpb_inst_8_dout[2]),
  .I1(sdpb_inst_9_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(sdpb_inst_10_dout[2]),
  .I1(sdpb_inst_11_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(sdpb_inst_12_dout[2]),
  .I1(sdpb_inst_13_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sdpb_inst_14_dout[2]),
  .I1(sdpb_inst_15_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(sdpb_inst_16_dout[2]),
  .I1(sdpb_inst_17_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(sdpb_inst_18_dout[2]),
  .I1(sdpb_inst_19_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(sdpb_inst_20_dout[2]),
  .I1(sdpb_inst_21_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(sdpb_inst_22_dout[2]),
  .I1(sdpb_inst_23_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(sdpb_inst_24_dout[2]),
  .I1(sdpb_inst_25_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(sdpb_inst_26_dout[2]),
  .I1(sdpb_inst_27_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(sdpb_inst_28_dout[2]),
  .I1(sdpb_inst_29_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(sdpb_inst_30_dout[2]),
  .I1(sdpb_inst_31_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(sdpb_inst_32_dout[2]),
  .I1(sdpb_inst_33_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(sdpb_inst_34_dout[2]),
  .I1(sdpb_inst_35_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(sdpb_inst_36_dout[2]),
  .I1(sdpb_inst_37_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(sdpb_inst_38_dout[2]),
  .I1(sdpb_inst_39_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(sdpb_inst_40_dout[2]),
  .I1(sdpb_inst_41_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(sdpb_inst_42_dout[2]),
  .I1(sdpb_inst_43_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(sdpb_inst_44_dout[2]),
  .I1(sdpb_inst_45_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(sdpb_inst_46_dout[2]),
  .I1(sdpb_inst_47_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(sdpb_inst_48_dout[2]),
  .I1(sdpb_inst_49_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(sdpb_inst_50_dout[2]),
  .I1(sdpb_inst_51_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(sdpb_inst_52_dout[2]),
  .I1(sdpb_inst_53_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(sdpb_inst_54_dout[2]),
  .I1(sdpb_inst_55_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(sdpb_inst_56_dout[2]),
  .I1(sdpb_inst_57_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(sdpb_inst_58_dout[2]),
  .I1(sdpb_inst_59_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(sdpb_inst_60_dout[2]),
  .I1(sdpb_inst_61_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(sdpb_inst_62_dout[2]),
  .I1(sdpb_inst_63_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(sdpb_inst_64_dout[2]),
  .I1(sdpb_inst_65_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(sdpb_inst_66_dout[2]),
  .I1(sdpb_inst_67_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(sdpb_inst_68_dout[2]),
  .I1(sdpb_inst_69_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(sdpb_inst_70_dout[2]),
  .I1(sdpb_inst_71_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(sdpb_inst_72_dout[2]),
  .I1(sdpb_inst_73_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(sdpb_inst_74_dout[2]),
  .I1(sdpb_inst_75_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(sdpb_inst_76_dout[2]),
  .I1(sdpb_inst_77_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(sdpb_inst_78_dout[2]),
  .I1(sdpb_inst_79_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(sdpb_inst_80_dout[2]),
  .I1(sdpb_inst_81_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(sdpb_inst_82_dout[2]),
  .I1(sdpb_inst_83_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(sdpb_inst_84_dout[2]),
  .I1(sdpb_inst_85_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(sdpb_inst_86_dout[2]),
  .I1(sdpb_inst_87_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(sdpb_inst_88_dout[2]),
  .I1(sdpb_inst_89_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(sdpb_inst_90_dout[2]),
  .I1(sdpb_inst_91_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(sdpb_inst_92_dout[2]),
  .I1(sdpb_inst_93_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(sdpb_inst_94_dout[2]),
  .I1(sdpb_inst_95_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(sdpb_inst_96_dout[2]),
  .I1(sdpb_inst_97_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(sdpb_inst_98_dout[2]),
  .I1(sdpb_inst_99_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(sdpb_inst_100_dout[2]),
  .I1(sdpb_inst_101_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(sdpb_inst_102_dout[2]),
  .I1(sdpb_inst_103_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(sdpb_inst_104_dout[2]),
  .I1(sdpb_inst_105_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(sdpb_inst_106_dout[2]),
  .I1(sdpb_inst_107_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(sdpb_inst_108_dout[2]),
  .I1(sdpb_inst_109_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(sdpb_inst_110_dout[2]),
  .I1(sdpb_inst_111_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(sdpb_inst_112_dout[2]),
  .I1(sdpb_inst_113_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(sdpb_inst_114_dout[2]),
  .I1(sdpb_inst_115_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(sdpb_inst_116_dout[2]),
  .I1(sdpb_inst_117_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(sdpb_inst_118_dout[2]),
  .I1(sdpb_inst_119_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(sdpb_inst_120_dout[2]),
  .I1(sdpb_inst_121_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sdpb_inst_122_dout[2]),
  .I1(sdpb_inst_123_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sdpb_inst_124_dout[2]),
  .I1(sdpb_inst_125_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sdpb_inst_126_dout[2]),
  .I1(sdpb_inst_127_dout[2]),
  .S0(dff_q_6)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_5)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_5)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(dff_q_5)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(dff_q_5)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(dff_q_5)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(dff_q_5)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_5)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_5)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_5)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_5)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_5)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_5)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(dff_q_5)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_5)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_5)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(dff_q_5)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_286),
  .I1(mux_o_287),
  .S0(dff_q_5)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(mux_o_288),
  .I1(mux_o_289),
  .S0(dff_q_5)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(mux_o_290),
  .I1(mux_o_291),
  .S0(dff_q_5)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(mux_o_292),
  .I1(mux_o_293),
  .S0(dff_q_5)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(dff_q_5)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(dff_q_5)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_5)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_5)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_5)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(dff_q_5)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(dff_q_5)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_5)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_5)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_5)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_314),
  .I1(mux_o_315),
  .S0(dff_q_5)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(dff_q_5)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_318),
  .I1(mux_o_319),
  .S0(dff_q_4)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(dff_q_4)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(dff_q_4)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(dff_q_4)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(dff_q_4)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_328),
  .I1(mux_o_329),
  .S0(dff_q_4)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(dff_q_4)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_4)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_4)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_4)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_4)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_4)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(dff_q_4)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(mux_o_344),
  .I1(mux_o_345),
  .S0(dff_q_4)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(mux_o_346),
  .I1(mux_o_347),
  .S0(dff_q_4)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(mux_o_348),
  .I1(mux_o_349),
  .S0(dff_q_4)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_3)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_3)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_3)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_356),
  .I1(mux_o_357),
  .S0(dff_q_3)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_358),
  .I1(mux_o_359),
  .S0(dff_q_3)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(dff_q_3)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_362),
  .I1(mux_o_363),
  .S0(dff_q_3)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_3)
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_2)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_2)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(dff_q_2)
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(dff_q_2)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(mux_o_374),
  .I1(mux_o_375),
  .S0(dff_q_1)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(mux_o_376),
  .I1(mux_o_377),
  .S0(dff_q_1)
);
MUX2 mux_inst_380 (
  .O(dout[2]),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(dff_q_0)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(sdpb_inst_0_dout[3]),
  .I1(sdpb_inst_1_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(sdpb_inst_2_dout[3]),
  .I1(sdpb_inst_3_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(sdpb_inst_4_dout[3]),
  .I1(sdpb_inst_5_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(sdpb_inst_6_dout[3]),
  .I1(sdpb_inst_7_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(sdpb_inst_8_dout[3]),
  .I1(sdpb_inst_9_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(sdpb_inst_10_dout[3]),
  .I1(sdpb_inst_11_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(sdpb_inst_12_dout[3]),
  .I1(sdpb_inst_13_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(sdpb_inst_14_dout[3]),
  .I1(sdpb_inst_15_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(sdpb_inst_16_dout[3]),
  .I1(sdpb_inst_17_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(sdpb_inst_18_dout[3]),
  .I1(sdpb_inst_19_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(sdpb_inst_20_dout[3]),
  .I1(sdpb_inst_21_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(sdpb_inst_22_dout[3]),
  .I1(sdpb_inst_23_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(sdpb_inst_24_dout[3]),
  .I1(sdpb_inst_25_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(sdpb_inst_26_dout[3]),
  .I1(sdpb_inst_27_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(sdpb_inst_28_dout[3]),
  .I1(sdpb_inst_29_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(sdpb_inst_30_dout[3]),
  .I1(sdpb_inst_31_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(sdpb_inst_32_dout[3]),
  .I1(sdpb_inst_33_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(sdpb_inst_34_dout[3]),
  .I1(sdpb_inst_35_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(sdpb_inst_36_dout[3]),
  .I1(sdpb_inst_37_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(sdpb_inst_38_dout[3]),
  .I1(sdpb_inst_39_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(sdpb_inst_40_dout[3]),
  .I1(sdpb_inst_41_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(sdpb_inst_42_dout[3]),
  .I1(sdpb_inst_43_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(sdpb_inst_44_dout[3]),
  .I1(sdpb_inst_45_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(sdpb_inst_46_dout[3]),
  .I1(sdpb_inst_47_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(sdpb_inst_48_dout[3]),
  .I1(sdpb_inst_49_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(sdpb_inst_50_dout[3]),
  .I1(sdpb_inst_51_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(sdpb_inst_52_dout[3]),
  .I1(sdpb_inst_53_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(sdpb_inst_54_dout[3]),
  .I1(sdpb_inst_55_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(sdpb_inst_56_dout[3]),
  .I1(sdpb_inst_57_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(sdpb_inst_58_dout[3]),
  .I1(sdpb_inst_59_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(sdpb_inst_60_dout[3]),
  .I1(sdpb_inst_61_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(sdpb_inst_62_dout[3]),
  .I1(sdpb_inst_63_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(sdpb_inst_64_dout[3]),
  .I1(sdpb_inst_65_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(sdpb_inst_66_dout[3]),
  .I1(sdpb_inst_67_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(sdpb_inst_68_dout[3]),
  .I1(sdpb_inst_69_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(sdpb_inst_70_dout[3]),
  .I1(sdpb_inst_71_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(sdpb_inst_72_dout[3]),
  .I1(sdpb_inst_73_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(sdpb_inst_74_dout[3]),
  .I1(sdpb_inst_75_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(sdpb_inst_76_dout[3]),
  .I1(sdpb_inst_77_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(sdpb_inst_78_dout[3]),
  .I1(sdpb_inst_79_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(sdpb_inst_80_dout[3]),
  .I1(sdpb_inst_81_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(sdpb_inst_82_dout[3]),
  .I1(sdpb_inst_83_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(sdpb_inst_84_dout[3]),
  .I1(sdpb_inst_85_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(sdpb_inst_86_dout[3]),
  .I1(sdpb_inst_87_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(sdpb_inst_88_dout[3]),
  .I1(sdpb_inst_89_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(sdpb_inst_90_dout[3]),
  .I1(sdpb_inst_91_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(sdpb_inst_92_dout[3]),
  .I1(sdpb_inst_93_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(sdpb_inst_94_dout[3]),
  .I1(sdpb_inst_95_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(sdpb_inst_96_dout[3]),
  .I1(sdpb_inst_97_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(sdpb_inst_98_dout[3]),
  .I1(sdpb_inst_99_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(sdpb_inst_100_dout[3]),
  .I1(sdpb_inst_101_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(sdpb_inst_102_dout[3]),
  .I1(sdpb_inst_103_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(sdpb_inst_104_dout[3]),
  .I1(sdpb_inst_105_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(sdpb_inst_106_dout[3]),
  .I1(sdpb_inst_107_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(sdpb_inst_108_dout[3]),
  .I1(sdpb_inst_109_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sdpb_inst_110_dout[3]),
  .I1(sdpb_inst_111_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(sdpb_inst_112_dout[3]),
  .I1(sdpb_inst_113_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(sdpb_inst_114_dout[3]),
  .I1(sdpb_inst_115_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(sdpb_inst_116_dout[3]),
  .I1(sdpb_inst_117_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sdpb_inst_118_dout[3]),
  .I1(sdpb_inst_119_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sdpb_inst_120_dout[3]),
  .I1(sdpb_inst_121_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sdpb_inst_122_dout[3]),
  .I1(sdpb_inst_123_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(sdpb_inst_124_dout[3]),
  .I1(sdpb_inst_125_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(sdpb_inst_126_dout[3]),
  .I1(sdpb_inst_127_dout[3]),
  .S0(dff_q_6)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_381),
  .I1(mux_o_382),
  .S0(dff_q_5)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_383),
  .I1(mux_o_384),
  .S0(dff_q_5)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_385),
  .I1(mux_o_386),
  .S0(dff_q_5)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(mux_o_387),
  .I1(mux_o_388),
  .S0(dff_q_5)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(mux_o_389),
  .I1(mux_o_390),
  .S0(dff_q_5)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(mux_o_391),
  .I1(mux_o_392),
  .S0(dff_q_5)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(mux_o_393),
  .I1(mux_o_394),
  .S0(dff_q_5)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(mux_o_395),
  .I1(mux_o_396),
  .S0(dff_q_5)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(mux_o_397),
  .I1(mux_o_398),
  .S0(dff_q_5)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_399),
  .I1(mux_o_400),
  .S0(dff_q_5)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_401),
  .I1(mux_o_402),
  .S0(dff_q_5)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_403),
  .I1(mux_o_404),
  .S0(dff_q_5)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(dff_q_5)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(dff_q_5)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_5)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(dff_q_5)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_5)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_5)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_5)
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(mux_o_419),
  .I1(mux_o_420),
  .S0(dff_q_5)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(mux_o_421),
  .I1(mux_o_422),
  .S0(dff_q_5)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(mux_o_423),
  .I1(mux_o_424),
  .S0(dff_q_5)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(mux_o_425),
  .I1(mux_o_426),
  .S0(dff_q_5)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(mux_o_427),
  .I1(mux_o_428),
  .S0(dff_q_5)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(mux_o_429),
  .I1(mux_o_430),
  .S0(dff_q_5)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(mux_o_431),
  .I1(mux_o_432),
  .S0(dff_q_5)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(mux_o_433),
  .I1(mux_o_434),
  .S0(dff_q_5)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(mux_o_435),
  .I1(mux_o_436),
  .S0(dff_q_5)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_437),
  .I1(mux_o_438),
  .S0(dff_q_5)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_439),
  .I1(mux_o_440),
  .S0(dff_q_5)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_5)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_5)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_4)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_4)
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(dff_q_4)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(dff_q_4)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_453),
  .I1(mux_o_454),
  .S0(dff_q_4)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_455),
  .I1(mux_o_456),
  .S0(dff_q_4)
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_457),
  .I1(mux_o_458),
  .S0(dff_q_4)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_459),
  .I1(mux_o_460),
  .S0(dff_q_4)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(dff_q_4)
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_463),
  .I1(mux_o_464),
  .S0(dff_q_4)
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_4)
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_4)
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_4)
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_4)
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_4)
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_4)
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_3)
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(dff_q_3)
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(dff_q_3)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(mux_o_483),
  .I1(mux_o_484),
  .S0(dff_q_3)
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(mux_o_485),
  .I1(mux_o_486),
  .S0(dff_q_3)
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(mux_o_487),
  .I1(mux_o_488),
  .S0(dff_q_3)
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(mux_o_489),
  .I1(mux_o_490),
  .S0(dff_q_3)
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(dff_q_3)
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(dff_q_2)
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(mux_o_495),
  .I1(mux_o_496),
  .S0(dff_q_2)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(mux_o_497),
  .I1(mux_o_498),
  .S0(dff_q_2)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(mux_o_499),
  .I1(mux_o_500),
  .S0(dff_q_2)
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(mux_o_501),
  .I1(mux_o_502),
  .S0(dff_q_1)
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(mux_o_503),
  .I1(mux_o_504),
  .S0(dff_q_1)
);
MUX2 mux_inst_507 (
  .O(dout[3]),
  .I0(mux_o_505),
  .I1(mux_o_506),
  .S0(dff_q_0)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(sdpb_inst_0_dout[4]),
  .I1(sdpb_inst_1_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(sdpb_inst_2_dout[4]),
  .I1(sdpb_inst_3_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(sdpb_inst_4_dout[4]),
  .I1(sdpb_inst_5_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(sdpb_inst_6_dout[4]),
  .I1(sdpb_inst_7_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(sdpb_inst_8_dout[4]),
  .I1(sdpb_inst_9_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(sdpb_inst_10_dout[4]),
  .I1(sdpb_inst_11_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(sdpb_inst_12_dout[4]),
  .I1(sdpb_inst_13_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(sdpb_inst_14_dout[4]),
  .I1(sdpb_inst_15_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(sdpb_inst_16_dout[4]),
  .I1(sdpb_inst_17_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(sdpb_inst_18_dout[4]),
  .I1(sdpb_inst_19_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(sdpb_inst_20_dout[4]),
  .I1(sdpb_inst_21_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(sdpb_inst_22_dout[4]),
  .I1(sdpb_inst_23_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(sdpb_inst_24_dout[4]),
  .I1(sdpb_inst_25_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(sdpb_inst_26_dout[4]),
  .I1(sdpb_inst_27_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(sdpb_inst_28_dout[4]),
  .I1(sdpb_inst_29_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(sdpb_inst_30_dout[4]),
  .I1(sdpb_inst_31_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(sdpb_inst_32_dout[4]),
  .I1(sdpb_inst_33_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(sdpb_inst_34_dout[4]),
  .I1(sdpb_inst_35_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(sdpb_inst_36_dout[4]),
  .I1(sdpb_inst_37_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(sdpb_inst_38_dout[4]),
  .I1(sdpb_inst_39_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(sdpb_inst_40_dout[4]),
  .I1(sdpb_inst_41_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(sdpb_inst_42_dout[4]),
  .I1(sdpb_inst_43_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(sdpb_inst_44_dout[4]),
  .I1(sdpb_inst_45_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(sdpb_inst_46_dout[4]),
  .I1(sdpb_inst_47_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(sdpb_inst_48_dout[4]),
  .I1(sdpb_inst_49_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(sdpb_inst_50_dout[4]),
  .I1(sdpb_inst_51_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(sdpb_inst_52_dout[4]),
  .I1(sdpb_inst_53_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(sdpb_inst_54_dout[4]),
  .I1(sdpb_inst_55_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(sdpb_inst_56_dout[4]),
  .I1(sdpb_inst_57_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(sdpb_inst_58_dout[4]),
  .I1(sdpb_inst_59_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(sdpb_inst_60_dout[4]),
  .I1(sdpb_inst_61_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(sdpb_inst_62_dout[4]),
  .I1(sdpb_inst_63_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(sdpb_inst_64_dout[4]),
  .I1(sdpb_inst_65_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(sdpb_inst_66_dout[4]),
  .I1(sdpb_inst_67_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(sdpb_inst_68_dout[4]),
  .I1(sdpb_inst_69_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(sdpb_inst_70_dout[4]),
  .I1(sdpb_inst_71_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(sdpb_inst_72_dout[4]),
  .I1(sdpb_inst_73_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(sdpb_inst_74_dout[4]),
  .I1(sdpb_inst_75_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(sdpb_inst_76_dout[4]),
  .I1(sdpb_inst_77_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(sdpb_inst_78_dout[4]),
  .I1(sdpb_inst_79_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(sdpb_inst_80_dout[4]),
  .I1(sdpb_inst_81_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(sdpb_inst_82_dout[4]),
  .I1(sdpb_inst_83_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(sdpb_inst_84_dout[4]),
  .I1(sdpb_inst_85_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(sdpb_inst_86_dout[4]),
  .I1(sdpb_inst_87_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(sdpb_inst_88_dout[4]),
  .I1(sdpb_inst_89_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(sdpb_inst_90_dout[4]),
  .I1(sdpb_inst_91_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(sdpb_inst_92_dout[4]),
  .I1(sdpb_inst_93_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(sdpb_inst_94_dout[4]),
  .I1(sdpb_inst_95_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(sdpb_inst_96_dout[4]),
  .I1(sdpb_inst_97_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(sdpb_inst_98_dout[4]),
  .I1(sdpb_inst_99_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(sdpb_inst_100_dout[4]),
  .I1(sdpb_inst_101_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(sdpb_inst_102_dout[4]),
  .I1(sdpb_inst_103_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(sdpb_inst_104_dout[4]),
  .I1(sdpb_inst_105_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(sdpb_inst_106_dout[4]),
  .I1(sdpb_inst_107_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(sdpb_inst_108_dout[4]),
  .I1(sdpb_inst_109_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(sdpb_inst_110_dout[4]),
  .I1(sdpb_inst_111_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(sdpb_inst_112_dout[4]),
  .I1(sdpb_inst_113_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(sdpb_inst_114_dout[4]),
  .I1(sdpb_inst_115_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(sdpb_inst_116_dout[4]),
  .I1(sdpb_inst_117_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(sdpb_inst_118_dout[4]),
  .I1(sdpb_inst_119_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(sdpb_inst_120_dout[4]),
  .I1(sdpb_inst_121_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(sdpb_inst_122_dout[4]),
  .I1(sdpb_inst_123_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(sdpb_inst_124_dout[4]),
  .I1(sdpb_inst_125_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(sdpb_inst_126_dout[4]),
  .I1(sdpb_inst_127_dout[4]),
  .S0(dff_q_6)
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(dff_q_5)
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(dff_q_5)
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(dff_q_5)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(dff_q_5)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(dff_q_5)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(dff_q_5)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(dff_q_5)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_5)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(dff_q_5)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_526),
  .I1(mux_o_527),
  .S0(dff_q_5)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_528),
  .I1(mux_o_529),
  .S0(dff_q_5)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_530),
  .I1(mux_o_531),
  .S0(dff_q_5)
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_532),
  .I1(mux_o_533),
  .S0(dff_q_5)
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(mux_o_534),
  .I1(mux_o_535),
  .S0(dff_q_5)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_536),
  .I1(mux_o_537),
  .S0(dff_q_5)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_538),
  .I1(mux_o_539),
  .S0(dff_q_5)
);
MUX2 mux_inst_588 (
  .O(mux_o_588),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(dff_q_5)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(mux_o_542),
  .I1(mux_o_543),
  .S0(dff_q_5)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(dff_q_5)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(mux_o_546),
  .I1(mux_o_547),
  .S0(dff_q_5)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(mux_o_548),
  .I1(mux_o_549),
  .S0(dff_q_5)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(mux_o_550),
  .I1(mux_o_551),
  .S0(dff_q_5)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(mux_o_552),
  .I1(mux_o_553),
  .S0(dff_q_5)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(mux_o_554),
  .I1(mux_o_555),
  .S0(dff_q_5)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(mux_o_556),
  .I1(mux_o_557),
  .S0(dff_q_5)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(dff_q_5)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(dff_q_5)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(dff_q_5)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(dff_q_5)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_566),
  .I1(mux_o_567),
  .S0(dff_q_5)
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(mux_o_568),
  .I1(mux_o_569),
  .S0(dff_q_5)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(mux_o_570),
  .I1(mux_o_571),
  .S0(dff_q_5)
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(dff_q_4)
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(dff_q_4)
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(dff_q_4)
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(dff_q_4)
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(dff_q_4)
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(dff_q_4)
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_584),
  .I1(mux_o_585),
  .S0(dff_q_4)
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(dff_q_4)
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_588),
  .I1(mux_o_589),
  .S0(dff_q_4)
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_590),
  .I1(mux_o_591),
  .S0(dff_q_4)
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_592),
  .I1(mux_o_593),
  .S0(dff_q_4)
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_594),
  .I1(mux_o_595),
  .S0(dff_q_4)
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_596),
  .I1(mux_o_597),
  .S0(dff_q_4)
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_598),
  .I1(mux_o_599),
  .S0(dff_q_4)
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_600),
  .I1(mux_o_601),
  .S0(dff_q_4)
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(mux_o_602),
  .I1(mux_o_603),
  .S0(dff_q_4)
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(mux_o_604),
  .I1(mux_o_605),
  .S0(dff_q_3)
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(mux_o_606),
  .I1(mux_o_607),
  .S0(dff_q_3)
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(mux_o_608),
  .I1(mux_o_609),
  .S0(dff_q_3)
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(mux_o_610),
  .I1(mux_o_611),
  .S0(dff_q_3)
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_612),
  .I1(mux_o_613),
  .S0(dff_q_3)
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_614),
  .I1(mux_o_615),
  .S0(dff_q_3)
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_616),
  .I1(mux_o_617),
  .S0(dff_q_3)
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(mux_o_618),
  .I1(mux_o_619),
  .S0(dff_q_3)
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_620),
  .I1(mux_o_621),
  .S0(dff_q_2)
);
MUX2 mux_inst_629 (
  .O(mux_o_629),
  .I0(mux_o_622),
  .I1(mux_o_623),
  .S0(dff_q_2)
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(mux_o_624),
  .I1(mux_o_625),
  .S0(dff_q_2)
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(mux_o_626),
  .I1(mux_o_627),
  .S0(dff_q_2)
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(mux_o_628),
  .I1(mux_o_629),
  .S0(dff_q_1)
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(dff_q_1)
);
MUX2 mux_inst_634 (
  .O(dout[4]),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(dff_q_0)
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(sdpb_inst_0_dout[5]),
  .I1(sdpb_inst_1_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(sdpb_inst_2_dout[5]),
  .I1(sdpb_inst_3_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(sdpb_inst_4_dout[5]),
  .I1(sdpb_inst_5_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(sdpb_inst_6_dout[5]),
  .I1(sdpb_inst_7_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(sdpb_inst_8_dout[5]),
  .I1(sdpb_inst_9_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(sdpb_inst_10_dout[5]),
  .I1(sdpb_inst_11_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(sdpb_inst_12_dout[5]),
  .I1(sdpb_inst_13_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(sdpb_inst_14_dout[5]),
  .I1(sdpb_inst_15_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(sdpb_inst_16_dout[5]),
  .I1(sdpb_inst_17_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(sdpb_inst_18_dout[5]),
  .I1(sdpb_inst_19_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(sdpb_inst_20_dout[5]),
  .I1(sdpb_inst_21_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(sdpb_inst_22_dout[5]),
  .I1(sdpb_inst_23_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(sdpb_inst_24_dout[5]),
  .I1(sdpb_inst_25_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(sdpb_inst_26_dout[5]),
  .I1(sdpb_inst_27_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(sdpb_inst_28_dout[5]),
  .I1(sdpb_inst_29_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(sdpb_inst_30_dout[5]),
  .I1(sdpb_inst_31_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(sdpb_inst_32_dout[5]),
  .I1(sdpb_inst_33_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(sdpb_inst_34_dout[5]),
  .I1(sdpb_inst_35_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(sdpb_inst_36_dout[5]),
  .I1(sdpb_inst_37_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(sdpb_inst_38_dout[5]),
  .I1(sdpb_inst_39_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(sdpb_inst_40_dout[5]),
  .I1(sdpb_inst_41_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(sdpb_inst_42_dout[5]),
  .I1(sdpb_inst_43_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(sdpb_inst_44_dout[5]),
  .I1(sdpb_inst_45_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(sdpb_inst_46_dout[5]),
  .I1(sdpb_inst_47_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(sdpb_inst_48_dout[5]),
  .I1(sdpb_inst_49_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(sdpb_inst_50_dout[5]),
  .I1(sdpb_inst_51_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(sdpb_inst_52_dout[5]),
  .I1(sdpb_inst_53_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(sdpb_inst_54_dout[5]),
  .I1(sdpb_inst_55_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(sdpb_inst_56_dout[5]),
  .I1(sdpb_inst_57_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(sdpb_inst_58_dout[5]),
  .I1(sdpb_inst_59_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(sdpb_inst_60_dout[5]),
  .I1(sdpb_inst_61_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(sdpb_inst_62_dout[5]),
  .I1(sdpb_inst_63_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(sdpb_inst_64_dout[5]),
  .I1(sdpb_inst_65_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(sdpb_inst_66_dout[5]),
  .I1(sdpb_inst_67_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(sdpb_inst_68_dout[5]),
  .I1(sdpb_inst_69_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(sdpb_inst_70_dout[5]),
  .I1(sdpb_inst_71_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(sdpb_inst_72_dout[5]),
  .I1(sdpb_inst_73_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(sdpb_inst_74_dout[5]),
  .I1(sdpb_inst_75_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(sdpb_inst_76_dout[5]),
  .I1(sdpb_inst_77_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(sdpb_inst_78_dout[5]),
  .I1(sdpb_inst_79_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(sdpb_inst_80_dout[5]),
  .I1(sdpb_inst_81_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(sdpb_inst_82_dout[5]),
  .I1(sdpb_inst_83_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(sdpb_inst_84_dout[5]),
  .I1(sdpb_inst_85_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(sdpb_inst_86_dout[5]),
  .I1(sdpb_inst_87_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(sdpb_inst_88_dout[5]),
  .I1(sdpb_inst_89_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(sdpb_inst_90_dout[5]),
  .I1(sdpb_inst_91_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(sdpb_inst_92_dout[5]),
  .I1(sdpb_inst_93_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(sdpb_inst_94_dout[5]),
  .I1(sdpb_inst_95_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(sdpb_inst_96_dout[5]),
  .I1(sdpb_inst_97_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(sdpb_inst_98_dout[5]),
  .I1(sdpb_inst_99_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(sdpb_inst_100_dout[5]),
  .I1(sdpb_inst_101_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(sdpb_inst_102_dout[5]),
  .I1(sdpb_inst_103_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(sdpb_inst_104_dout[5]),
  .I1(sdpb_inst_105_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(sdpb_inst_106_dout[5]),
  .I1(sdpb_inst_107_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(sdpb_inst_108_dout[5]),
  .I1(sdpb_inst_109_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(sdpb_inst_110_dout[5]),
  .I1(sdpb_inst_111_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(sdpb_inst_112_dout[5]),
  .I1(sdpb_inst_113_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(sdpb_inst_114_dout[5]),
  .I1(sdpb_inst_115_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(sdpb_inst_116_dout[5]),
  .I1(sdpb_inst_117_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(sdpb_inst_118_dout[5]),
  .I1(sdpb_inst_119_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(sdpb_inst_120_dout[5]),
  .I1(sdpb_inst_121_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(sdpb_inst_122_dout[5]),
  .I1(sdpb_inst_123_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(sdpb_inst_124_dout[5]),
  .I1(sdpb_inst_125_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(sdpb_inst_126_dout[5]),
  .I1(sdpb_inst_127_dout[5]),
  .S0(dff_q_6)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_635),
  .I1(mux_o_636),
  .S0(dff_q_5)
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_637),
  .I1(mux_o_638),
  .S0(dff_q_5)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_639),
  .I1(mux_o_640),
  .S0(dff_q_5)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_641),
  .I1(mux_o_642),
  .S0(dff_q_5)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_643),
  .I1(mux_o_644),
  .S0(dff_q_5)
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(mux_o_645),
  .I1(mux_o_646),
  .S0(dff_q_5)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(mux_o_647),
  .I1(mux_o_648),
  .S0(dff_q_5)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(mux_o_649),
  .I1(mux_o_650),
  .S0(dff_q_5)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(mux_o_651),
  .I1(mux_o_652),
  .S0(dff_q_5)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_653),
  .I1(mux_o_654),
  .S0(dff_q_5)
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(mux_o_655),
  .I1(mux_o_656),
  .S0(dff_q_5)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(mux_o_657),
  .I1(mux_o_658),
  .S0(dff_q_5)
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(mux_o_659),
  .I1(mux_o_660),
  .S0(dff_q_5)
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(mux_o_661),
  .I1(mux_o_662),
  .S0(dff_q_5)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(mux_o_663),
  .I1(mux_o_664),
  .S0(dff_q_5)
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(mux_o_665),
  .I1(mux_o_666),
  .S0(dff_q_5)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(mux_o_667),
  .I1(mux_o_668),
  .S0(dff_q_5)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(mux_o_669),
  .I1(mux_o_670),
  .S0(dff_q_5)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(mux_o_671),
  .I1(mux_o_672),
  .S0(dff_q_5)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(mux_o_673),
  .I1(mux_o_674),
  .S0(dff_q_5)
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(mux_o_675),
  .I1(mux_o_676),
  .S0(dff_q_5)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(mux_o_677),
  .I1(mux_o_678),
  .S0(dff_q_5)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(mux_o_679),
  .I1(mux_o_680),
  .S0(dff_q_5)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(mux_o_681),
  .I1(mux_o_682),
  .S0(dff_q_5)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(mux_o_683),
  .I1(mux_o_684),
  .S0(dff_q_5)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(mux_o_685),
  .I1(mux_o_686),
  .S0(dff_q_5)
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(mux_o_687),
  .I1(mux_o_688),
  .S0(dff_q_5)
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(mux_o_689),
  .I1(mux_o_690),
  .S0(dff_q_5)
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(mux_o_691),
  .I1(mux_o_692),
  .S0(dff_q_5)
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(mux_o_693),
  .I1(mux_o_694),
  .S0(dff_q_5)
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_695),
  .I1(mux_o_696),
  .S0(dff_q_5)
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_697),
  .I1(mux_o_698),
  .S0(dff_q_5)
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_699),
  .I1(mux_o_700),
  .S0(dff_q_4)
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_701),
  .I1(mux_o_702),
  .S0(dff_q_4)
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_703),
  .I1(mux_o_704),
  .S0(dff_q_4)
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(dff_q_4)
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_707),
  .I1(mux_o_708),
  .S0(dff_q_4)
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_709),
  .I1(mux_o_710),
  .S0(dff_q_4)
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_711),
  .I1(mux_o_712),
  .S0(dff_q_4)
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(dff_q_4)
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_4)
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_4)
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(dff_q_4)
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(dff_q_4)
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(dff_q_4)
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(mux_o_725),
  .I1(mux_o_726),
  .S0(dff_q_4)
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(mux_o_727),
  .I1(mux_o_728),
  .S0(dff_q_4)
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(dff_q_4)
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(dff_q_3)
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(dff_q_3)
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(dff_q_3)
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(dff_q_3)
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(dff_q_3)
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(dff_q_3)
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(mux_o_743),
  .I1(mux_o_744),
  .S0(dff_q_3)
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(mux_o_745),
  .I1(mux_o_746),
  .S0(dff_q_3)
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(mux_o_747),
  .I1(mux_o_748),
  .S0(dff_q_2)
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(mux_o_749),
  .I1(mux_o_750),
  .S0(dff_q_2)
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(mux_o_751),
  .I1(mux_o_752),
  .S0(dff_q_2)
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(mux_o_753),
  .I1(mux_o_754),
  .S0(dff_q_2)
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(mux_o_755),
  .I1(mux_o_756),
  .S0(dff_q_1)
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(mux_o_757),
  .I1(mux_o_758),
  .S0(dff_q_1)
);
MUX2 mux_inst_761 (
  .O(dout[5]),
  .I0(mux_o_759),
  .I1(mux_o_760),
  .S0(dff_q_0)
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(sdpb_inst_0_dout[6]),
  .I1(sdpb_inst_1_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(sdpb_inst_2_dout[6]),
  .I1(sdpb_inst_3_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(sdpb_inst_4_dout[6]),
  .I1(sdpb_inst_5_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(sdpb_inst_6_dout[6]),
  .I1(sdpb_inst_7_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(sdpb_inst_8_dout[6]),
  .I1(sdpb_inst_9_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(sdpb_inst_10_dout[6]),
  .I1(sdpb_inst_11_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(sdpb_inst_12_dout[6]),
  .I1(sdpb_inst_13_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(sdpb_inst_14_dout[6]),
  .I1(sdpb_inst_15_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(sdpb_inst_16_dout[6]),
  .I1(sdpb_inst_17_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(sdpb_inst_18_dout[6]),
  .I1(sdpb_inst_19_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(sdpb_inst_20_dout[6]),
  .I1(sdpb_inst_21_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(sdpb_inst_22_dout[6]),
  .I1(sdpb_inst_23_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(sdpb_inst_24_dout[6]),
  .I1(sdpb_inst_25_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(sdpb_inst_26_dout[6]),
  .I1(sdpb_inst_27_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(sdpb_inst_28_dout[6]),
  .I1(sdpb_inst_29_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(sdpb_inst_30_dout[6]),
  .I1(sdpb_inst_31_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(sdpb_inst_32_dout[6]),
  .I1(sdpb_inst_33_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(sdpb_inst_34_dout[6]),
  .I1(sdpb_inst_35_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(sdpb_inst_36_dout[6]),
  .I1(sdpb_inst_37_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(sdpb_inst_38_dout[6]),
  .I1(sdpb_inst_39_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(sdpb_inst_40_dout[6]),
  .I1(sdpb_inst_41_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(sdpb_inst_42_dout[6]),
  .I1(sdpb_inst_43_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(sdpb_inst_44_dout[6]),
  .I1(sdpb_inst_45_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(sdpb_inst_46_dout[6]),
  .I1(sdpb_inst_47_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(sdpb_inst_48_dout[6]),
  .I1(sdpb_inst_49_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(sdpb_inst_50_dout[6]),
  .I1(sdpb_inst_51_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(sdpb_inst_52_dout[6]),
  .I1(sdpb_inst_53_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(sdpb_inst_54_dout[6]),
  .I1(sdpb_inst_55_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(sdpb_inst_56_dout[6]),
  .I1(sdpb_inst_57_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(sdpb_inst_58_dout[6]),
  .I1(sdpb_inst_59_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(sdpb_inst_60_dout[6]),
  .I1(sdpb_inst_61_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(sdpb_inst_62_dout[6]),
  .I1(sdpb_inst_63_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(sdpb_inst_64_dout[6]),
  .I1(sdpb_inst_65_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(sdpb_inst_66_dout[6]),
  .I1(sdpb_inst_67_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(sdpb_inst_68_dout[6]),
  .I1(sdpb_inst_69_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(sdpb_inst_70_dout[6]),
  .I1(sdpb_inst_71_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(sdpb_inst_72_dout[6]),
  .I1(sdpb_inst_73_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(sdpb_inst_74_dout[6]),
  .I1(sdpb_inst_75_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(sdpb_inst_76_dout[6]),
  .I1(sdpb_inst_77_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(sdpb_inst_78_dout[6]),
  .I1(sdpb_inst_79_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(sdpb_inst_80_dout[6]),
  .I1(sdpb_inst_81_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(sdpb_inst_82_dout[6]),
  .I1(sdpb_inst_83_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(sdpb_inst_84_dout[6]),
  .I1(sdpb_inst_85_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(sdpb_inst_86_dout[6]),
  .I1(sdpb_inst_87_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(sdpb_inst_88_dout[6]),
  .I1(sdpb_inst_89_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(sdpb_inst_90_dout[6]),
  .I1(sdpb_inst_91_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(sdpb_inst_92_dout[6]),
  .I1(sdpb_inst_93_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(sdpb_inst_94_dout[6]),
  .I1(sdpb_inst_95_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(sdpb_inst_96_dout[6]),
  .I1(sdpb_inst_97_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(sdpb_inst_98_dout[6]),
  .I1(sdpb_inst_99_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(sdpb_inst_100_dout[6]),
  .I1(sdpb_inst_101_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(sdpb_inst_102_dout[6]),
  .I1(sdpb_inst_103_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(sdpb_inst_104_dout[6]),
  .I1(sdpb_inst_105_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(sdpb_inst_106_dout[6]),
  .I1(sdpb_inst_107_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(sdpb_inst_108_dout[6]),
  .I1(sdpb_inst_109_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(sdpb_inst_110_dout[6]),
  .I1(sdpb_inst_111_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(sdpb_inst_112_dout[6]),
  .I1(sdpb_inst_113_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(sdpb_inst_114_dout[6]),
  .I1(sdpb_inst_115_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(sdpb_inst_116_dout[6]),
  .I1(sdpb_inst_117_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(sdpb_inst_118_dout[6]),
  .I1(sdpb_inst_119_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(sdpb_inst_120_dout[6]),
  .I1(sdpb_inst_121_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(sdpb_inst_122_dout[6]),
  .I1(sdpb_inst_123_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(sdpb_inst_124_dout[6]),
  .I1(sdpb_inst_125_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(sdpb_inst_126_dout[6]),
  .I1(sdpb_inst_127_dout[6]),
  .S0(dff_q_6)
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(dff_q_5)
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(dff_q_5)
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(dff_q_5)
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(dff_q_5)
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(dff_q_5)
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(dff_q_5)
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(mux_o_774),
  .I1(mux_o_775),
  .S0(dff_q_5)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(mux_o_776),
  .I1(mux_o_777),
  .S0(dff_q_5)
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(mux_o_778),
  .I1(mux_o_779),
  .S0(dff_q_5)
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(mux_o_780),
  .I1(mux_o_781),
  .S0(dff_q_5)
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(mux_o_782),
  .I1(mux_o_783),
  .S0(dff_q_5)
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(mux_o_784),
  .I1(mux_o_785),
  .S0(dff_q_5)
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(mux_o_786),
  .I1(mux_o_787),
  .S0(dff_q_5)
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(mux_o_788),
  .I1(mux_o_789),
  .S0(dff_q_5)
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(mux_o_790),
  .I1(mux_o_791),
  .S0(dff_q_5)
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(dff_q_5)
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(mux_o_794),
  .I1(mux_o_795),
  .S0(dff_q_5)
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(mux_o_796),
  .I1(mux_o_797),
  .S0(dff_q_5)
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(mux_o_798),
  .I1(mux_o_799),
  .S0(dff_q_5)
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(mux_o_800),
  .I1(mux_o_801),
  .S0(dff_q_5)
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(mux_o_802),
  .I1(mux_o_803),
  .S0(dff_q_5)
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(mux_o_804),
  .I1(mux_o_805),
  .S0(dff_q_5)
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(dff_q_5)
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(dff_q_5)
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(dff_q_5)
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(dff_q_5)
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(dff_q_5)
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(dff_q_5)
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(dff_q_5)
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(dff_q_5)
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(dff_q_5)
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(mux_o_824),
  .I1(mux_o_825),
  .S0(dff_q_5)
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(mux_o_826),
  .I1(mux_o_827),
  .S0(dff_q_4)
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(mux_o_828),
  .I1(mux_o_829),
  .S0(dff_q_4)
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(mux_o_830),
  .I1(mux_o_831),
  .S0(dff_q_4)
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(mux_o_832),
  .I1(mux_o_833),
  .S0(dff_q_4)
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(mux_o_834),
  .I1(mux_o_835),
  .S0(dff_q_4)
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_836),
  .I1(mux_o_837),
  .S0(dff_q_4)
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_838),
  .I1(mux_o_839),
  .S0(dff_q_4)
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_840),
  .I1(mux_o_841),
  .S0(dff_q_4)
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_842),
  .I1(mux_o_843),
  .S0(dff_q_4)
);
MUX2 mux_inst_867 (
  .O(mux_o_867),
  .I0(mux_o_844),
  .I1(mux_o_845),
  .S0(dff_q_4)
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(mux_o_846),
  .I1(mux_o_847),
  .S0(dff_q_4)
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(mux_o_848),
  .I1(mux_o_849),
  .S0(dff_q_4)
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(mux_o_850),
  .I1(mux_o_851),
  .S0(dff_q_4)
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(mux_o_852),
  .I1(mux_o_853),
  .S0(dff_q_4)
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(mux_o_854),
  .I1(mux_o_855),
  .S0(dff_q_4)
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(mux_o_856),
  .I1(mux_o_857),
  .S0(dff_q_4)
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(mux_o_858),
  .I1(mux_o_859),
  .S0(dff_q_3)
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(mux_o_860),
  .I1(mux_o_861),
  .S0(dff_q_3)
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(mux_o_862),
  .I1(mux_o_863),
  .S0(dff_q_3)
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(mux_o_864),
  .I1(mux_o_865),
  .S0(dff_q_3)
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(mux_o_866),
  .I1(mux_o_867),
  .S0(dff_q_3)
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(mux_o_868),
  .I1(mux_o_869),
  .S0(dff_q_3)
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(mux_o_870),
  .I1(mux_o_871),
  .S0(dff_q_3)
);
MUX2 mux_inst_881 (
  .O(mux_o_881),
  .I0(mux_o_872),
  .I1(mux_o_873),
  .S0(dff_q_3)
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(mux_o_874),
  .I1(mux_o_875),
  .S0(dff_q_2)
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(mux_o_876),
  .I1(mux_o_877),
  .S0(dff_q_2)
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(mux_o_878),
  .I1(mux_o_879),
  .S0(dff_q_2)
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(mux_o_880),
  .I1(mux_o_881),
  .S0(dff_q_2)
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(dff_q_1)
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(dff_q_1)
);
MUX2 mux_inst_888 (
  .O(dout[6]),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(dff_q_0)
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(sdpb_inst_0_dout[7]),
  .I1(sdpb_inst_1_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(sdpb_inst_2_dout[7]),
  .I1(sdpb_inst_3_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(sdpb_inst_4_dout[7]),
  .I1(sdpb_inst_5_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(sdpb_inst_6_dout[7]),
  .I1(sdpb_inst_7_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(sdpb_inst_8_dout[7]),
  .I1(sdpb_inst_9_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(sdpb_inst_10_dout[7]),
  .I1(sdpb_inst_11_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(sdpb_inst_12_dout[7]),
  .I1(sdpb_inst_13_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(sdpb_inst_14_dout[7]),
  .I1(sdpb_inst_15_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(sdpb_inst_16_dout[7]),
  .I1(sdpb_inst_17_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_898 (
  .O(mux_o_898),
  .I0(sdpb_inst_18_dout[7]),
  .I1(sdpb_inst_19_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(sdpb_inst_20_dout[7]),
  .I1(sdpb_inst_21_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(sdpb_inst_22_dout[7]),
  .I1(sdpb_inst_23_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(sdpb_inst_24_dout[7]),
  .I1(sdpb_inst_25_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(sdpb_inst_26_dout[7]),
  .I1(sdpb_inst_27_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(sdpb_inst_28_dout[7]),
  .I1(sdpb_inst_29_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(sdpb_inst_30_dout[7]),
  .I1(sdpb_inst_31_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(sdpb_inst_32_dout[7]),
  .I1(sdpb_inst_33_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(sdpb_inst_34_dout[7]),
  .I1(sdpb_inst_35_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(sdpb_inst_36_dout[7]),
  .I1(sdpb_inst_37_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(sdpb_inst_38_dout[7]),
  .I1(sdpb_inst_39_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(sdpb_inst_40_dout[7]),
  .I1(sdpb_inst_41_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(sdpb_inst_42_dout[7]),
  .I1(sdpb_inst_43_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(sdpb_inst_44_dout[7]),
  .I1(sdpb_inst_45_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(sdpb_inst_46_dout[7]),
  .I1(sdpb_inst_47_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(sdpb_inst_48_dout[7]),
  .I1(sdpb_inst_49_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(sdpb_inst_50_dout[7]),
  .I1(sdpb_inst_51_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(sdpb_inst_52_dout[7]),
  .I1(sdpb_inst_53_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(sdpb_inst_54_dout[7]),
  .I1(sdpb_inst_55_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(sdpb_inst_56_dout[7]),
  .I1(sdpb_inst_57_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(sdpb_inst_58_dout[7]),
  .I1(sdpb_inst_59_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(sdpb_inst_60_dout[7]),
  .I1(sdpb_inst_61_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(sdpb_inst_62_dout[7]),
  .I1(sdpb_inst_63_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(sdpb_inst_64_dout[7]),
  .I1(sdpb_inst_65_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(sdpb_inst_66_dout[7]),
  .I1(sdpb_inst_67_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(sdpb_inst_68_dout[7]),
  .I1(sdpb_inst_69_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(sdpb_inst_70_dout[7]),
  .I1(sdpb_inst_71_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(sdpb_inst_72_dout[7]),
  .I1(sdpb_inst_73_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(sdpb_inst_74_dout[7]),
  .I1(sdpb_inst_75_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(sdpb_inst_76_dout[7]),
  .I1(sdpb_inst_77_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(sdpb_inst_78_dout[7]),
  .I1(sdpb_inst_79_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_929 (
  .O(mux_o_929),
  .I0(sdpb_inst_80_dout[7]),
  .I1(sdpb_inst_81_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(sdpb_inst_82_dout[7]),
  .I1(sdpb_inst_83_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(sdpb_inst_84_dout[7]),
  .I1(sdpb_inst_85_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(sdpb_inst_86_dout[7]),
  .I1(sdpb_inst_87_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(sdpb_inst_88_dout[7]),
  .I1(sdpb_inst_89_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(sdpb_inst_90_dout[7]),
  .I1(sdpb_inst_91_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(sdpb_inst_92_dout[7]),
  .I1(sdpb_inst_93_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(sdpb_inst_94_dout[7]),
  .I1(sdpb_inst_95_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(sdpb_inst_96_dout[7]),
  .I1(sdpb_inst_97_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(sdpb_inst_98_dout[7]),
  .I1(sdpb_inst_99_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(sdpb_inst_100_dout[7]),
  .I1(sdpb_inst_101_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(sdpb_inst_102_dout[7]),
  .I1(sdpb_inst_103_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(sdpb_inst_104_dout[7]),
  .I1(sdpb_inst_105_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(sdpb_inst_106_dout[7]),
  .I1(sdpb_inst_107_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(sdpb_inst_108_dout[7]),
  .I1(sdpb_inst_109_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_944 (
  .O(mux_o_944),
  .I0(sdpb_inst_110_dout[7]),
  .I1(sdpb_inst_111_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(sdpb_inst_112_dout[7]),
  .I1(sdpb_inst_113_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(sdpb_inst_114_dout[7]),
  .I1(sdpb_inst_115_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(sdpb_inst_116_dout[7]),
  .I1(sdpb_inst_117_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(sdpb_inst_118_dout[7]),
  .I1(sdpb_inst_119_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(sdpb_inst_120_dout[7]),
  .I1(sdpb_inst_121_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(sdpb_inst_122_dout[7]),
  .I1(sdpb_inst_123_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(sdpb_inst_124_dout[7]),
  .I1(sdpb_inst_125_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(sdpb_inst_126_dout[7]),
  .I1(sdpb_inst_127_dout[7]),
  .S0(dff_q_6)
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(mux_o_889),
  .I1(mux_o_890),
  .S0(dff_q_5)
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(mux_o_891),
  .I1(mux_o_892),
  .S0(dff_q_5)
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(mux_o_893),
  .I1(mux_o_894),
  .S0(dff_q_5)
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(mux_o_895),
  .I1(mux_o_896),
  .S0(dff_q_5)
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(mux_o_897),
  .I1(mux_o_898),
  .S0(dff_q_5)
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(mux_o_899),
  .I1(mux_o_900),
  .S0(dff_q_5)
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(mux_o_901),
  .I1(mux_o_902),
  .S0(dff_q_5)
);
MUX2 mux_inst_960 (
  .O(mux_o_960),
  .I0(mux_o_903),
  .I1(mux_o_904),
  .S0(dff_q_5)
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(mux_o_905),
  .I1(mux_o_906),
  .S0(dff_q_5)
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(mux_o_907),
  .I1(mux_o_908),
  .S0(dff_q_5)
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(mux_o_909),
  .I1(mux_o_910),
  .S0(dff_q_5)
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(mux_o_911),
  .I1(mux_o_912),
  .S0(dff_q_5)
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(mux_o_913),
  .I1(mux_o_914),
  .S0(dff_q_5)
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(mux_o_915),
  .I1(mux_o_916),
  .S0(dff_q_5)
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(mux_o_917),
  .I1(mux_o_918),
  .S0(dff_q_5)
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(mux_o_919),
  .I1(mux_o_920),
  .S0(dff_q_5)
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(mux_o_921),
  .I1(mux_o_922),
  .S0(dff_q_5)
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(mux_o_923),
  .I1(mux_o_924),
  .S0(dff_q_5)
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(mux_o_925),
  .I1(mux_o_926),
  .S0(dff_q_5)
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(mux_o_927),
  .I1(mux_o_928),
  .S0(dff_q_5)
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(mux_o_929),
  .I1(mux_o_930),
  .S0(dff_q_5)
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(mux_o_931),
  .I1(mux_o_932),
  .S0(dff_q_5)
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(mux_o_933),
  .I1(mux_o_934),
  .S0(dff_q_5)
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(mux_o_935),
  .I1(mux_o_936),
  .S0(dff_q_5)
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(mux_o_937),
  .I1(mux_o_938),
  .S0(dff_q_5)
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(mux_o_939),
  .I1(mux_o_940),
  .S0(dff_q_5)
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(mux_o_941),
  .I1(mux_o_942),
  .S0(dff_q_5)
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(mux_o_943),
  .I1(mux_o_944),
  .S0(dff_q_5)
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(mux_o_945),
  .I1(mux_o_946),
  .S0(dff_q_5)
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(mux_o_947),
  .I1(mux_o_948),
  .S0(dff_q_5)
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(mux_o_949),
  .I1(mux_o_950),
  .S0(dff_q_5)
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(mux_o_951),
  .I1(mux_o_952),
  .S0(dff_q_5)
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(mux_o_953),
  .I1(mux_o_954),
  .S0(dff_q_4)
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(mux_o_955),
  .I1(mux_o_956),
  .S0(dff_q_4)
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(mux_o_957),
  .I1(mux_o_958),
  .S0(dff_q_4)
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(mux_o_959),
  .I1(mux_o_960),
  .S0(dff_q_4)
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(dff_q_4)
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(dff_q_4)
);
MUX2 mux_inst_991 (
  .O(mux_o_991),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(dff_q_4)
);
MUX2 mux_inst_992 (
  .O(mux_o_992),
  .I0(mux_o_967),
  .I1(mux_o_968),
  .S0(dff_q_4)
);
MUX2 mux_inst_993 (
  .O(mux_o_993),
  .I0(mux_o_969),
  .I1(mux_o_970),
  .S0(dff_q_4)
);
MUX2 mux_inst_994 (
  .O(mux_o_994),
  .I0(mux_o_971),
  .I1(mux_o_972),
  .S0(dff_q_4)
);
MUX2 mux_inst_995 (
  .O(mux_o_995),
  .I0(mux_o_973),
  .I1(mux_o_974),
  .S0(dff_q_4)
);
MUX2 mux_inst_996 (
  .O(mux_o_996),
  .I0(mux_o_975),
  .I1(mux_o_976),
  .S0(dff_q_4)
);
MUX2 mux_inst_997 (
  .O(mux_o_997),
  .I0(mux_o_977),
  .I1(mux_o_978),
  .S0(dff_q_4)
);
MUX2 mux_inst_998 (
  .O(mux_o_998),
  .I0(mux_o_979),
  .I1(mux_o_980),
  .S0(dff_q_4)
);
MUX2 mux_inst_999 (
  .O(mux_o_999),
  .I0(mux_o_981),
  .I1(mux_o_982),
  .S0(dff_q_4)
);
MUX2 mux_inst_1000 (
  .O(mux_o_1000),
  .I0(mux_o_983),
  .I1(mux_o_984),
  .S0(dff_q_4)
);
MUX2 mux_inst_1001 (
  .O(mux_o_1001),
  .I0(mux_o_985),
  .I1(mux_o_986),
  .S0(dff_q_3)
);
MUX2 mux_inst_1002 (
  .O(mux_o_1002),
  .I0(mux_o_987),
  .I1(mux_o_988),
  .S0(dff_q_3)
);
MUX2 mux_inst_1003 (
  .O(mux_o_1003),
  .I0(mux_o_989),
  .I1(mux_o_990),
  .S0(dff_q_3)
);
MUX2 mux_inst_1004 (
  .O(mux_o_1004),
  .I0(mux_o_991),
  .I1(mux_o_992),
  .S0(dff_q_3)
);
MUX2 mux_inst_1005 (
  .O(mux_o_1005),
  .I0(mux_o_993),
  .I1(mux_o_994),
  .S0(dff_q_3)
);
MUX2 mux_inst_1006 (
  .O(mux_o_1006),
  .I0(mux_o_995),
  .I1(mux_o_996),
  .S0(dff_q_3)
);
MUX2 mux_inst_1007 (
  .O(mux_o_1007),
  .I0(mux_o_997),
  .I1(mux_o_998),
  .S0(dff_q_3)
);
MUX2 mux_inst_1008 (
  .O(mux_o_1008),
  .I0(mux_o_999),
  .I1(mux_o_1000),
  .S0(dff_q_3)
);
MUX2 mux_inst_1009 (
  .O(mux_o_1009),
  .I0(mux_o_1001),
  .I1(mux_o_1002),
  .S0(dff_q_2)
);
MUX2 mux_inst_1010 (
  .O(mux_o_1010),
  .I0(mux_o_1003),
  .I1(mux_o_1004),
  .S0(dff_q_2)
);
MUX2 mux_inst_1011 (
  .O(mux_o_1011),
  .I0(mux_o_1005),
  .I1(mux_o_1006),
  .S0(dff_q_2)
);
MUX2 mux_inst_1012 (
  .O(mux_o_1012),
  .I0(mux_o_1007),
  .I1(mux_o_1008),
  .S0(dff_q_2)
);
MUX2 mux_inst_1013 (
  .O(mux_o_1013),
  .I0(mux_o_1009),
  .I1(mux_o_1010),
  .S0(dff_q_1)
);
MUX2 mux_inst_1014 (
  .O(mux_o_1014),
  .I0(mux_o_1011),
  .I1(mux_o_1012),
  .S0(dff_q_1)
);
MUX2 mux_inst_1015 (
  .O(dout[7]),
  .I0(mux_o_1013),
  .I1(mux_o_1014),
  .S0(dff_q_0)
);
MUX2 mux_inst_1016 (
  .O(mux_o_1016),
  .I0(sdpb_inst_0_dout[8]),
  .I1(sdpb_inst_1_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1017 (
  .O(mux_o_1017),
  .I0(sdpb_inst_2_dout[8]),
  .I1(sdpb_inst_3_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1018 (
  .O(mux_o_1018),
  .I0(sdpb_inst_4_dout[8]),
  .I1(sdpb_inst_5_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1019 (
  .O(mux_o_1019),
  .I0(sdpb_inst_6_dout[8]),
  .I1(sdpb_inst_7_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1020 (
  .O(mux_o_1020),
  .I0(sdpb_inst_8_dout[8]),
  .I1(sdpb_inst_9_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1021 (
  .O(mux_o_1021),
  .I0(sdpb_inst_10_dout[8]),
  .I1(sdpb_inst_11_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1022 (
  .O(mux_o_1022),
  .I0(sdpb_inst_12_dout[8]),
  .I1(sdpb_inst_13_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1023 (
  .O(mux_o_1023),
  .I0(sdpb_inst_14_dout[8]),
  .I1(sdpb_inst_15_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1024 (
  .O(mux_o_1024),
  .I0(sdpb_inst_16_dout[8]),
  .I1(sdpb_inst_17_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1025 (
  .O(mux_o_1025),
  .I0(sdpb_inst_18_dout[8]),
  .I1(sdpb_inst_19_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1026 (
  .O(mux_o_1026),
  .I0(sdpb_inst_20_dout[8]),
  .I1(sdpb_inst_21_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1027 (
  .O(mux_o_1027),
  .I0(sdpb_inst_22_dout[8]),
  .I1(sdpb_inst_23_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1028 (
  .O(mux_o_1028),
  .I0(sdpb_inst_24_dout[8]),
  .I1(sdpb_inst_25_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1029 (
  .O(mux_o_1029),
  .I0(sdpb_inst_26_dout[8]),
  .I1(sdpb_inst_27_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1030 (
  .O(mux_o_1030),
  .I0(sdpb_inst_28_dout[8]),
  .I1(sdpb_inst_29_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1031 (
  .O(mux_o_1031),
  .I0(sdpb_inst_30_dout[8]),
  .I1(sdpb_inst_31_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1032 (
  .O(mux_o_1032),
  .I0(sdpb_inst_32_dout[8]),
  .I1(sdpb_inst_33_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1033 (
  .O(mux_o_1033),
  .I0(sdpb_inst_34_dout[8]),
  .I1(sdpb_inst_35_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1034 (
  .O(mux_o_1034),
  .I0(sdpb_inst_36_dout[8]),
  .I1(sdpb_inst_37_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1035 (
  .O(mux_o_1035),
  .I0(sdpb_inst_38_dout[8]),
  .I1(sdpb_inst_39_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1036 (
  .O(mux_o_1036),
  .I0(sdpb_inst_40_dout[8]),
  .I1(sdpb_inst_41_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1037 (
  .O(mux_o_1037),
  .I0(sdpb_inst_42_dout[8]),
  .I1(sdpb_inst_43_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1038 (
  .O(mux_o_1038),
  .I0(sdpb_inst_44_dout[8]),
  .I1(sdpb_inst_45_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1039 (
  .O(mux_o_1039),
  .I0(sdpb_inst_46_dout[8]),
  .I1(sdpb_inst_47_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1040 (
  .O(mux_o_1040),
  .I0(sdpb_inst_48_dout[8]),
  .I1(sdpb_inst_49_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1041 (
  .O(mux_o_1041),
  .I0(sdpb_inst_50_dout[8]),
  .I1(sdpb_inst_51_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1042 (
  .O(mux_o_1042),
  .I0(sdpb_inst_52_dout[8]),
  .I1(sdpb_inst_53_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1043 (
  .O(mux_o_1043),
  .I0(sdpb_inst_54_dout[8]),
  .I1(sdpb_inst_55_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1044 (
  .O(mux_o_1044),
  .I0(sdpb_inst_56_dout[8]),
  .I1(sdpb_inst_57_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1045 (
  .O(mux_o_1045),
  .I0(sdpb_inst_58_dout[8]),
  .I1(sdpb_inst_59_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1046 (
  .O(mux_o_1046),
  .I0(sdpb_inst_60_dout[8]),
  .I1(sdpb_inst_61_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1047 (
  .O(mux_o_1047),
  .I0(sdpb_inst_62_dout[8]),
  .I1(sdpb_inst_63_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1048 (
  .O(mux_o_1048),
  .I0(sdpb_inst_64_dout[8]),
  .I1(sdpb_inst_65_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1049 (
  .O(mux_o_1049),
  .I0(sdpb_inst_66_dout[8]),
  .I1(sdpb_inst_67_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1050 (
  .O(mux_o_1050),
  .I0(sdpb_inst_68_dout[8]),
  .I1(sdpb_inst_69_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1051 (
  .O(mux_o_1051),
  .I0(sdpb_inst_70_dout[8]),
  .I1(sdpb_inst_71_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1052 (
  .O(mux_o_1052),
  .I0(sdpb_inst_72_dout[8]),
  .I1(sdpb_inst_73_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1053 (
  .O(mux_o_1053),
  .I0(sdpb_inst_74_dout[8]),
  .I1(sdpb_inst_75_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1054 (
  .O(mux_o_1054),
  .I0(sdpb_inst_76_dout[8]),
  .I1(sdpb_inst_77_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1055 (
  .O(mux_o_1055),
  .I0(sdpb_inst_78_dout[8]),
  .I1(sdpb_inst_79_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1056 (
  .O(mux_o_1056),
  .I0(sdpb_inst_80_dout[8]),
  .I1(sdpb_inst_81_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1057 (
  .O(mux_o_1057),
  .I0(sdpb_inst_82_dout[8]),
  .I1(sdpb_inst_83_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1058 (
  .O(mux_o_1058),
  .I0(sdpb_inst_84_dout[8]),
  .I1(sdpb_inst_85_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1059 (
  .O(mux_o_1059),
  .I0(sdpb_inst_86_dout[8]),
  .I1(sdpb_inst_87_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1060 (
  .O(mux_o_1060),
  .I0(sdpb_inst_88_dout[8]),
  .I1(sdpb_inst_89_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1061 (
  .O(mux_o_1061),
  .I0(sdpb_inst_90_dout[8]),
  .I1(sdpb_inst_91_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1062 (
  .O(mux_o_1062),
  .I0(sdpb_inst_92_dout[8]),
  .I1(sdpb_inst_93_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1063 (
  .O(mux_o_1063),
  .I0(sdpb_inst_94_dout[8]),
  .I1(sdpb_inst_95_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1064 (
  .O(mux_o_1064),
  .I0(sdpb_inst_96_dout[8]),
  .I1(sdpb_inst_97_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1065 (
  .O(mux_o_1065),
  .I0(sdpb_inst_98_dout[8]),
  .I1(sdpb_inst_99_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1066 (
  .O(mux_o_1066),
  .I0(sdpb_inst_100_dout[8]),
  .I1(sdpb_inst_101_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1067 (
  .O(mux_o_1067),
  .I0(sdpb_inst_102_dout[8]),
  .I1(sdpb_inst_103_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1068 (
  .O(mux_o_1068),
  .I0(sdpb_inst_104_dout[8]),
  .I1(sdpb_inst_105_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1069 (
  .O(mux_o_1069),
  .I0(sdpb_inst_106_dout[8]),
  .I1(sdpb_inst_107_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1070 (
  .O(mux_o_1070),
  .I0(sdpb_inst_108_dout[8]),
  .I1(sdpb_inst_109_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1071 (
  .O(mux_o_1071),
  .I0(sdpb_inst_110_dout[8]),
  .I1(sdpb_inst_111_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1072 (
  .O(mux_o_1072),
  .I0(sdpb_inst_112_dout[8]),
  .I1(sdpb_inst_113_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1073 (
  .O(mux_o_1073),
  .I0(sdpb_inst_114_dout[8]),
  .I1(sdpb_inst_115_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1074 (
  .O(mux_o_1074),
  .I0(sdpb_inst_116_dout[8]),
  .I1(sdpb_inst_117_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1075 (
  .O(mux_o_1075),
  .I0(sdpb_inst_118_dout[8]),
  .I1(sdpb_inst_119_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1076 (
  .O(mux_o_1076),
  .I0(sdpb_inst_120_dout[8]),
  .I1(sdpb_inst_121_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1077 (
  .O(mux_o_1077),
  .I0(sdpb_inst_122_dout[8]),
  .I1(sdpb_inst_123_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1078 (
  .O(mux_o_1078),
  .I0(sdpb_inst_124_dout[8]),
  .I1(sdpb_inst_125_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1079 (
  .O(mux_o_1079),
  .I0(sdpb_inst_126_dout[8]),
  .I1(sdpb_inst_127_dout[8]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1080 (
  .O(mux_o_1080),
  .I0(mux_o_1016),
  .I1(mux_o_1017),
  .S0(dff_q_5)
);
MUX2 mux_inst_1081 (
  .O(mux_o_1081),
  .I0(mux_o_1018),
  .I1(mux_o_1019),
  .S0(dff_q_5)
);
MUX2 mux_inst_1082 (
  .O(mux_o_1082),
  .I0(mux_o_1020),
  .I1(mux_o_1021),
  .S0(dff_q_5)
);
MUX2 mux_inst_1083 (
  .O(mux_o_1083),
  .I0(mux_o_1022),
  .I1(mux_o_1023),
  .S0(dff_q_5)
);
MUX2 mux_inst_1084 (
  .O(mux_o_1084),
  .I0(mux_o_1024),
  .I1(mux_o_1025),
  .S0(dff_q_5)
);
MUX2 mux_inst_1085 (
  .O(mux_o_1085),
  .I0(mux_o_1026),
  .I1(mux_o_1027),
  .S0(dff_q_5)
);
MUX2 mux_inst_1086 (
  .O(mux_o_1086),
  .I0(mux_o_1028),
  .I1(mux_o_1029),
  .S0(dff_q_5)
);
MUX2 mux_inst_1087 (
  .O(mux_o_1087),
  .I0(mux_o_1030),
  .I1(mux_o_1031),
  .S0(dff_q_5)
);
MUX2 mux_inst_1088 (
  .O(mux_o_1088),
  .I0(mux_o_1032),
  .I1(mux_o_1033),
  .S0(dff_q_5)
);
MUX2 mux_inst_1089 (
  .O(mux_o_1089),
  .I0(mux_o_1034),
  .I1(mux_o_1035),
  .S0(dff_q_5)
);
MUX2 mux_inst_1090 (
  .O(mux_o_1090),
  .I0(mux_o_1036),
  .I1(mux_o_1037),
  .S0(dff_q_5)
);
MUX2 mux_inst_1091 (
  .O(mux_o_1091),
  .I0(mux_o_1038),
  .I1(mux_o_1039),
  .S0(dff_q_5)
);
MUX2 mux_inst_1092 (
  .O(mux_o_1092),
  .I0(mux_o_1040),
  .I1(mux_o_1041),
  .S0(dff_q_5)
);
MUX2 mux_inst_1093 (
  .O(mux_o_1093),
  .I0(mux_o_1042),
  .I1(mux_o_1043),
  .S0(dff_q_5)
);
MUX2 mux_inst_1094 (
  .O(mux_o_1094),
  .I0(mux_o_1044),
  .I1(mux_o_1045),
  .S0(dff_q_5)
);
MUX2 mux_inst_1095 (
  .O(mux_o_1095),
  .I0(mux_o_1046),
  .I1(mux_o_1047),
  .S0(dff_q_5)
);
MUX2 mux_inst_1096 (
  .O(mux_o_1096),
  .I0(mux_o_1048),
  .I1(mux_o_1049),
  .S0(dff_q_5)
);
MUX2 mux_inst_1097 (
  .O(mux_o_1097),
  .I0(mux_o_1050),
  .I1(mux_o_1051),
  .S0(dff_q_5)
);
MUX2 mux_inst_1098 (
  .O(mux_o_1098),
  .I0(mux_o_1052),
  .I1(mux_o_1053),
  .S0(dff_q_5)
);
MUX2 mux_inst_1099 (
  .O(mux_o_1099),
  .I0(mux_o_1054),
  .I1(mux_o_1055),
  .S0(dff_q_5)
);
MUX2 mux_inst_1100 (
  .O(mux_o_1100),
  .I0(mux_o_1056),
  .I1(mux_o_1057),
  .S0(dff_q_5)
);
MUX2 mux_inst_1101 (
  .O(mux_o_1101),
  .I0(mux_o_1058),
  .I1(mux_o_1059),
  .S0(dff_q_5)
);
MUX2 mux_inst_1102 (
  .O(mux_o_1102),
  .I0(mux_o_1060),
  .I1(mux_o_1061),
  .S0(dff_q_5)
);
MUX2 mux_inst_1103 (
  .O(mux_o_1103),
  .I0(mux_o_1062),
  .I1(mux_o_1063),
  .S0(dff_q_5)
);
MUX2 mux_inst_1104 (
  .O(mux_o_1104),
  .I0(mux_o_1064),
  .I1(mux_o_1065),
  .S0(dff_q_5)
);
MUX2 mux_inst_1105 (
  .O(mux_o_1105),
  .I0(mux_o_1066),
  .I1(mux_o_1067),
  .S0(dff_q_5)
);
MUX2 mux_inst_1106 (
  .O(mux_o_1106),
  .I0(mux_o_1068),
  .I1(mux_o_1069),
  .S0(dff_q_5)
);
MUX2 mux_inst_1107 (
  .O(mux_o_1107),
  .I0(mux_o_1070),
  .I1(mux_o_1071),
  .S0(dff_q_5)
);
MUX2 mux_inst_1108 (
  .O(mux_o_1108),
  .I0(mux_o_1072),
  .I1(mux_o_1073),
  .S0(dff_q_5)
);
MUX2 mux_inst_1109 (
  .O(mux_o_1109),
  .I0(mux_o_1074),
  .I1(mux_o_1075),
  .S0(dff_q_5)
);
MUX2 mux_inst_1110 (
  .O(mux_o_1110),
  .I0(mux_o_1076),
  .I1(mux_o_1077),
  .S0(dff_q_5)
);
MUX2 mux_inst_1111 (
  .O(mux_o_1111),
  .I0(mux_o_1078),
  .I1(mux_o_1079),
  .S0(dff_q_5)
);
MUX2 mux_inst_1112 (
  .O(mux_o_1112),
  .I0(mux_o_1080),
  .I1(mux_o_1081),
  .S0(dff_q_4)
);
MUX2 mux_inst_1113 (
  .O(mux_o_1113),
  .I0(mux_o_1082),
  .I1(mux_o_1083),
  .S0(dff_q_4)
);
MUX2 mux_inst_1114 (
  .O(mux_o_1114),
  .I0(mux_o_1084),
  .I1(mux_o_1085),
  .S0(dff_q_4)
);
MUX2 mux_inst_1115 (
  .O(mux_o_1115),
  .I0(mux_o_1086),
  .I1(mux_o_1087),
  .S0(dff_q_4)
);
MUX2 mux_inst_1116 (
  .O(mux_o_1116),
  .I0(mux_o_1088),
  .I1(mux_o_1089),
  .S0(dff_q_4)
);
MUX2 mux_inst_1117 (
  .O(mux_o_1117),
  .I0(mux_o_1090),
  .I1(mux_o_1091),
  .S0(dff_q_4)
);
MUX2 mux_inst_1118 (
  .O(mux_o_1118),
  .I0(mux_o_1092),
  .I1(mux_o_1093),
  .S0(dff_q_4)
);
MUX2 mux_inst_1119 (
  .O(mux_o_1119),
  .I0(mux_o_1094),
  .I1(mux_o_1095),
  .S0(dff_q_4)
);
MUX2 mux_inst_1120 (
  .O(mux_o_1120),
  .I0(mux_o_1096),
  .I1(mux_o_1097),
  .S0(dff_q_4)
);
MUX2 mux_inst_1121 (
  .O(mux_o_1121),
  .I0(mux_o_1098),
  .I1(mux_o_1099),
  .S0(dff_q_4)
);
MUX2 mux_inst_1122 (
  .O(mux_o_1122),
  .I0(mux_o_1100),
  .I1(mux_o_1101),
  .S0(dff_q_4)
);
MUX2 mux_inst_1123 (
  .O(mux_o_1123),
  .I0(mux_o_1102),
  .I1(mux_o_1103),
  .S0(dff_q_4)
);
MUX2 mux_inst_1124 (
  .O(mux_o_1124),
  .I0(mux_o_1104),
  .I1(mux_o_1105),
  .S0(dff_q_4)
);
MUX2 mux_inst_1125 (
  .O(mux_o_1125),
  .I0(mux_o_1106),
  .I1(mux_o_1107),
  .S0(dff_q_4)
);
MUX2 mux_inst_1126 (
  .O(mux_o_1126),
  .I0(mux_o_1108),
  .I1(mux_o_1109),
  .S0(dff_q_4)
);
MUX2 mux_inst_1127 (
  .O(mux_o_1127),
  .I0(mux_o_1110),
  .I1(mux_o_1111),
  .S0(dff_q_4)
);
MUX2 mux_inst_1128 (
  .O(mux_o_1128),
  .I0(mux_o_1112),
  .I1(mux_o_1113),
  .S0(dff_q_3)
);
MUX2 mux_inst_1129 (
  .O(mux_o_1129),
  .I0(mux_o_1114),
  .I1(mux_o_1115),
  .S0(dff_q_3)
);
MUX2 mux_inst_1130 (
  .O(mux_o_1130),
  .I0(mux_o_1116),
  .I1(mux_o_1117),
  .S0(dff_q_3)
);
MUX2 mux_inst_1131 (
  .O(mux_o_1131),
  .I0(mux_o_1118),
  .I1(mux_o_1119),
  .S0(dff_q_3)
);
MUX2 mux_inst_1132 (
  .O(mux_o_1132),
  .I0(mux_o_1120),
  .I1(mux_o_1121),
  .S0(dff_q_3)
);
MUX2 mux_inst_1133 (
  .O(mux_o_1133),
  .I0(mux_o_1122),
  .I1(mux_o_1123),
  .S0(dff_q_3)
);
MUX2 mux_inst_1134 (
  .O(mux_o_1134),
  .I0(mux_o_1124),
  .I1(mux_o_1125),
  .S0(dff_q_3)
);
MUX2 mux_inst_1135 (
  .O(mux_o_1135),
  .I0(mux_o_1126),
  .I1(mux_o_1127),
  .S0(dff_q_3)
);
MUX2 mux_inst_1136 (
  .O(mux_o_1136),
  .I0(mux_o_1128),
  .I1(mux_o_1129),
  .S0(dff_q_2)
);
MUX2 mux_inst_1137 (
  .O(mux_o_1137),
  .I0(mux_o_1130),
  .I1(mux_o_1131),
  .S0(dff_q_2)
);
MUX2 mux_inst_1138 (
  .O(mux_o_1138),
  .I0(mux_o_1132),
  .I1(mux_o_1133),
  .S0(dff_q_2)
);
MUX2 mux_inst_1139 (
  .O(mux_o_1139),
  .I0(mux_o_1134),
  .I1(mux_o_1135),
  .S0(dff_q_2)
);
MUX2 mux_inst_1140 (
  .O(mux_o_1140),
  .I0(mux_o_1136),
  .I1(mux_o_1137),
  .S0(dff_q_1)
);
MUX2 mux_inst_1141 (
  .O(mux_o_1141),
  .I0(mux_o_1138),
  .I1(mux_o_1139),
  .S0(dff_q_1)
);
MUX2 mux_inst_1142 (
  .O(dout[8]),
  .I0(mux_o_1140),
  .I1(mux_o_1141),
  .S0(dff_q_0)
);
MUX2 mux_inst_1143 (
  .O(mux_o_1143),
  .I0(sdpb_inst_0_dout[9]),
  .I1(sdpb_inst_1_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1144 (
  .O(mux_o_1144),
  .I0(sdpb_inst_2_dout[9]),
  .I1(sdpb_inst_3_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1145 (
  .O(mux_o_1145),
  .I0(sdpb_inst_4_dout[9]),
  .I1(sdpb_inst_5_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1146 (
  .O(mux_o_1146),
  .I0(sdpb_inst_6_dout[9]),
  .I1(sdpb_inst_7_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1147 (
  .O(mux_o_1147),
  .I0(sdpb_inst_8_dout[9]),
  .I1(sdpb_inst_9_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1148 (
  .O(mux_o_1148),
  .I0(sdpb_inst_10_dout[9]),
  .I1(sdpb_inst_11_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1149 (
  .O(mux_o_1149),
  .I0(sdpb_inst_12_dout[9]),
  .I1(sdpb_inst_13_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1150 (
  .O(mux_o_1150),
  .I0(sdpb_inst_14_dout[9]),
  .I1(sdpb_inst_15_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1151 (
  .O(mux_o_1151),
  .I0(sdpb_inst_16_dout[9]),
  .I1(sdpb_inst_17_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1152 (
  .O(mux_o_1152),
  .I0(sdpb_inst_18_dout[9]),
  .I1(sdpb_inst_19_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1153 (
  .O(mux_o_1153),
  .I0(sdpb_inst_20_dout[9]),
  .I1(sdpb_inst_21_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1154 (
  .O(mux_o_1154),
  .I0(sdpb_inst_22_dout[9]),
  .I1(sdpb_inst_23_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1155 (
  .O(mux_o_1155),
  .I0(sdpb_inst_24_dout[9]),
  .I1(sdpb_inst_25_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1156 (
  .O(mux_o_1156),
  .I0(sdpb_inst_26_dout[9]),
  .I1(sdpb_inst_27_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1157 (
  .O(mux_o_1157),
  .I0(sdpb_inst_28_dout[9]),
  .I1(sdpb_inst_29_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1158 (
  .O(mux_o_1158),
  .I0(sdpb_inst_30_dout[9]),
  .I1(sdpb_inst_31_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1159 (
  .O(mux_o_1159),
  .I0(sdpb_inst_32_dout[9]),
  .I1(sdpb_inst_33_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1160 (
  .O(mux_o_1160),
  .I0(sdpb_inst_34_dout[9]),
  .I1(sdpb_inst_35_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1161 (
  .O(mux_o_1161),
  .I0(sdpb_inst_36_dout[9]),
  .I1(sdpb_inst_37_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1162 (
  .O(mux_o_1162),
  .I0(sdpb_inst_38_dout[9]),
  .I1(sdpb_inst_39_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1163 (
  .O(mux_o_1163),
  .I0(sdpb_inst_40_dout[9]),
  .I1(sdpb_inst_41_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1164 (
  .O(mux_o_1164),
  .I0(sdpb_inst_42_dout[9]),
  .I1(sdpb_inst_43_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1165 (
  .O(mux_o_1165),
  .I0(sdpb_inst_44_dout[9]),
  .I1(sdpb_inst_45_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1166 (
  .O(mux_o_1166),
  .I0(sdpb_inst_46_dout[9]),
  .I1(sdpb_inst_47_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1167 (
  .O(mux_o_1167),
  .I0(sdpb_inst_48_dout[9]),
  .I1(sdpb_inst_49_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1168 (
  .O(mux_o_1168),
  .I0(sdpb_inst_50_dout[9]),
  .I1(sdpb_inst_51_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1169 (
  .O(mux_o_1169),
  .I0(sdpb_inst_52_dout[9]),
  .I1(sdpb_inst_53_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1170 (
  .O(mux_o_1170),
  .I0(sdpb_inst_54_dout[9]),
  .I1(sdpb_inst_55_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1171 (
  .O(mux_o_1171),
  .I0(sdpb_inst_56_dout[9]),
  .I1(sdpb_inst_57_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1172 (
  .O(mux_o_1172),
  .I0(sdpb_inst_58_dout[9]),
  .I1(sdpb_inst_59_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1173 (
  .O(mux_o_1173),
  .I0(sdpb_inst_60_dout[9]),
  .I1(sdpb_inst_61_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1174 (
  .O(mux_o_1174),
  .I0(sdpb_inst_62_dout[9]),
  .I1(sdpb_inst_63_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1175 (
  .O(mux_o_1175),
  .I0(sdpb_inst_64_dout[9]),
  .I1(sdpb_inst_65_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1176 (
  .O(mux_o_1176),
  .I0(sdpb_inst_66_dout[9]),
  .I1(sdpb_inst_67_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1177 (
  .O(mux_o_1177),
  .I0(sdpb_inst_68_dout[9]),
  .I1(sdpb_inst_69_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1178 (
  .O(mux_o_1178),
  .I0(sdpb_inst_70_dout[9]),
  .I1(sdpb_inst_71_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1179 (
  .O(mux_o_1179),
  .I0(sdpb_inst_72_dout[9]),
  .I1(sdpb_inst_73_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1180 (
  .O(mux_o_1180),
  .I0(sdpb_inst_74_dout[9]),
  .I1(sdpb_inst_75_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1181 (
  .O(mux_o_1181),
  .I0(sdpb_inst_76_dout[9]),
  .I1(sdpb_inst_77_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1182 (
  .O(mux_o_1182),
  .I0(sdpb_inst_78_dout[9]),
  .I1(sdpb_inst_79_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1183 (
  .O(mux_o_1183),
  .I0(sdpb_inst_80_dout[9]),
  .I1(sdpb_inst_81_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1184 (
  .O(mux_o_1184),
  .I0(sdpb_inst_82_dout[9]),
  .I1(sdpb_inst_83_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1185 (
  .O(mux_o_1185),
  .I0(sdpb_inst_84_dout[9]),
  .I1(sdpb_inst_85_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1186 (
  .O(mux_o_1186),
  .I0(sdpb_inst_86_dout[9]),
  .I1(sdpb_inst_87_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1187 (
  .O(mux_o_1187),
  .I0(sdpb_inst_88_dout[9]),
  .I1(sdpb_inst_89_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1188 (
  .O(mux_o_1188),
  .I0(sdpb_inst_90_dout[9]),
  .I1(sdpb_inst_91_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1189 (
  .O(mux_o_1189),
  .I0(sdpb_inst_92_dout[9]),
  .I1(sdpb_inst_93_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1190 (
  .O(mux_o_1190),
  .I0(sdpb_inst_94_dout[9]),
  .I1(sdpb_inst_95_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1191 (
  .O(mux_o_1191),
  .I0(sdpb_inst_96_dout[9]),
  .I1(sdpb_inst_97_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1192 (
  .O(mux_o_1192),
  .I0(sdpb_inst_98_dout[9]),
  .I1(sdpb_inst_99_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1193 (
  .O(mux_o_1193),
  .I0(sdpb_inst_100_dout[9]),
  .I1(sdpb_inst_101_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1194 (
  .O(mux_o_1194),
  .I0(sdpb_inst_102_dout[9]),
  .I1(sdpb_inst_103_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1195 (
  .O(mux_o_1195),
  .I0(sdpb_inst_104_dout[9]),
  .I1(sdpb_inst_105_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1196 (
  .O(mux_o_1196),
  .I0(sdpb_inst_106_dout[9]),
  .I1(sdpb_inst_107_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1197 (
  .O(mux_o_1197),
  .I0(sdpb_inst_108_dout[9]),
  .I1(sdpb_inst_109_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1198 (
  .O(mux_o_1198),
  .I0(sdpb_inst_110_dout[9]),
  .I1(sdpb_inst_111_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1199 (
  .O(mux_o_1199),
  .I0(sdpb_inst_112_dout[9]),
  .I1(sdpb_inst_113_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1200 (
  .O(mux_o_1200),
  .I0(sdpb_inst_114_dout[9]),
  .I1(sdpb_inst_115_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1201 (
  .O(mux_o_1201),
  .I0(sdpb_inst_116_dout[9]),
  .I1(sdpb_inst_117_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1202 (
  .O(mux_o_1202),
  .I0(sdpb_inst_118_dout[9]),
  .I1(sdpb_inst_119_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1203 (
  .O(mux_o_1203),
  .I0(sdpb_inst_120_dout[9]),
  .I1(sdpb_inst_121_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1204 (
  .O(mux_o_1204),
  .I0(sdpb_inst_122_dout[9]),
  .I1(sdpb_inst_123_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1205 (
  .O(mux_o_1205),
  .I0(sdpb_inst_124_dout[9]),
  .I1(sdpb_inst_125_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1206 (
  .O(mux_o_1206),
  .I0(sdpb_inst_126_dout[9]),
  .I1(sdpb_inst_127_dout[9]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1207 (
  .O(mux_o_1207),
  .I0(mux_o_1143),
  .I1(mux_o_1144),
  .S0(dff_q_5)
);
MUX2 mux_inst_1208 (
  .O(mux_o_1208),
  .I0(mux_o_1145),
  .I1(mux_o_1146),
  .S0(dff_q_5)
);
MUX2 mux_inst_1209 (
  .O(mux_o_1209),
  .I0(mux_o_1147),
  .I1(mux_o_1148),
  .S0(dff_q_5)
);
MUX2 mux_inst_1210 (
  .O(mux_o_1210),
  .I0(mux_o_1149),
  .I1(mux_o_1150),
  .S0(dff_q_5)
);
MUX2 mux_inst_1211 (
  .O(mux_o_1211),
  .I0(mux_o_1151),
  .I1(mux_o_1152),
  .S0(dff_q_5)
);
MUX2 mux_inst_1212 (
  .O(mux_o_1212),
  .I0(mux_o_1153),
  .I1(mux_o_1154),
  .S0(dff_q_5)
);
MUX2 mux_inst_1213 (
  .O(mux_o_1213),
  .I0(mux_o_1155),
  .I1(mux_o_1156),
  .S0(dff_q_5)
);
MUX2 mux_inst_1214 (
  .O(mux_o_1214),
  .I0(mux_o_1157),
  .I1(mux_o_1158),
  .S0(dff_q_5)
);
MUX2 mux_inst_1215 (
  .O(mux_o_1215),
  .I0(mux_o_1159),
  .I1(mux_o_1160),
  .S0(dff_q_5)
);
MUX2 mux_inst_1216 (
  .O(mux_o_1216),
  .I0(mux_o_1161),
  .I1(mux_o_1162),
  .S0(dff_q_5)
);
MUX2 mux_inst_1217 (
  .O(mux_o_1217),
  .I0(mux_o_1163),
  .I1(mux_o_1164),
  .S0(dff_q_5)
);
MUX2 mux_inst_1218 (
  .O(mux_o_1218),
  .I0(mux_o_1165),
  .I1(mux_o_1166),
  .S0(dff_q_5)
);
MUX2 mux_inst_1219 (
  .O(mux_o_1219),
  .I0(mux_o_1167),
  .I1(mux_o_1168),
  .S0(dff_q_5)
);
MUX2 mux_inst_1220 (
  .O(mux_o_1220),
  .I0(mux_o_1169),
  .I1(mux_o_1170),
  .S0(dff_q_5)
);
MUX2 mux_inst_1221 (
  .O(mux_o_1221),
  .I0(mux_o_1171),
  .I1(mux_o_1172),
  .S0(dff_q_5)
);
MUX2 mux_inst_1222 (
  .O(mux_o_1222),
  .I0(mux_o_1173),
  .I1(mux_o_1174),
  .S0(dff_q_5)
);
MUX2 mux_inst_1223 (
  .O(mux_o_1223),
  .I0(mux_o_1175),
  .I1(mux_o_1176),
  .S0(dff_q_5)
);
MUX2 mux_inst_1224 (
  .O(mux_o_1224),
  .I0(mux_o_1177),
  .I1(mux_o_1178),
  .S0(dff_q_5)
);
MUX2 mux_inst_1225 (
  .O(mux_o_1225),
  .I0(mux_o_1179),
  .I1(mux_o_1180),
  .S0(dff_q_5)
);
MUX2 mux_inst_1226 (
  .O(mux_o_1226),
  .I0(mux_o_1181),
  .I1(mux_o_1182),
  .S0(dff_q_5)
);
MUX2 mux_inst_1227 (
  .O(mux_o_1227),
  .I0(mux_o_1183),
  .I1(mux_o_1184),
  .S0(dff_q_5)
);
MUX2 mux_inst_1228 (
  .O(mux_o_1228),
  .I0(mux_o_1185),
  .I1(mux_o_1186),
  .S0(dff_q_5)
);
MUX2 mux_inst_1229 (
  .O(mux_o_1229),
  .I0(mux_o_1187),
  .I1(mux_o_1188),
  .S0(dff_q_5)
);
MUX2 mux_inst_1230 (
  .O(mux_o_1230),
  .I0(mux_o_1189),
  .I1(mux_o_1190),
  .S0(dff_q_5)
);
MUX2 mux_inst_1231 (
  .O(mux_o_1231),
  .I0(mux_o_1191),
  .I1(mux_o_1192),
  .S0(dff_q_5)
);
MUX2 mux_inst_1232 (
  .O(mux_o_1232),
  .I0(mux_o_1193),
  .I1(mux_o_1194),
  .S0(dff_q_5)
);
MUX2 mux_inst_1233 (
  .O(mux_o_1233),
  .I0(mux_o_1195),
  .I1(mux_o_1196),
  .S0(dff_q_5)
);
MUX2 mux_inst_1234 (
  .O(mux_o_1234),
  .I0(mux_o_1197),
  .I1(mux_o_1198),
  .S0(dff_q_5)
);
MUX2 mux_inst_1235 (
  .O(mux_o_1235),
  .I0(mux_o_1199),
  .I1(mux_o_1200),
  .S0(dff_q_5)
);
MUX2 mux_inst_1236 (
  .O(mux_o_1236),
  .I0(mux_o_1201),
  .I1(mux_o_1202),
  .S0(dff_q_5)
);
MUX2 mux_inst_1237 (
  .O(mux_o_1237),
  .I0(mux_o_1203),
  .I1(mux_o_1204),
  .S0(dff_q_5)
);
MUX2 mux_inst_1238 (
  .O(mux_o_1238),
  .I0(mux_o_1205),
  .I1(mux_o_1206),
  .S0(dff_q_5)
);
MUX2 mux_inst_1239 (
  .O(mux_o_1239),
  .I0(mux_o_1207),
  .I1(mux_o_1208),
  .S0(dff_q_4)
);
MUX2 mux_inst_1240 (
  .O(mux_o_1240),
  .I0(mux_o_1209),
  .I1(mux_o_1210),
  .S0(dff_q_4)
);
MUX2 mux_inst_1241 (
  .O(mux_o_1241),
  .I0(mux_o_1211),
  .I1(mux_o_1212),
  .S0(dff_q_4)
);
MUX2 mux_inst_1242 (
  .O(mux_o_1242),
  .I0(mux_o_1213),
  .I1(mux_o_1214),
  .S0(dff_q_4)
);
MUX2 mux_inst_1243 (
  .O(mux_o_1243),
  .I0(mux_o_1215),
  .I1(mux_o_1216),
  .S0(dff_q_4)
);
MUX2 mux_inst_1244 (
  .O(mux_o_1244),
  .I0(mux_o_1217),
  .I1(mux_o_1218),
  .S0(dff_q_4)
);
MUX2 mux_inst_1245 (
  .O(mux_o_1245),
  .I0(mux_o_1219),
  .I1(mux_o_1220),
  .S0(dff_q_4)
);
MUX2 mux_inst_1246 (
  .O(mux_o_1246),
  .I0(mux_o_1221),
  .I1(mux_o_1222),
  .S0(dff_q_4)
);
MUX2 mux_inst_1247 (
  .O(mux_o_1247),
  .I0(mux_o_1223),
  .I1(mux_o_1224),
  .S0(dff_q_4)
);
MUX2 mux_inst_1248 (
  .O(mux_o_1248),
  .I0(mux_o_1225),
  .I1(mux_o_1226),
  .S0(dff_q_4)
);
MUX2 mux_inst_1249 (
  .O(mux_o_1249),
  .I0(mux_o_1227),
  .I1(mux_o_1228),
  .S0(dff_q_4)
);
MUX2 mux_inst_1250 (
  .O(mux_o_1250),
  .I0(mux_o_1229),
  .I1(mux_o_1230),
  .S0(dff_q_4)
);
MUX2 mux_inst_1251 (
  .O(mux_o_1251),
  .I0(mux_o_1231),
  .I1(mux_o_1232),
  .S0(dff_q_4)
);
MUX2 mux_inst_1252 (
  .O(mux_o_1252),
  .I0(mux_o_1233),
  .I1(mux_o_1234),
  .S0(dff_q_4)
);
MUX2 mux_inst_1253 (
  .O(mux_o_1253),
  .I0(mux_o_1235),
  .I1(mux_o_1236),
  .S0(dff_q_4)
);
MUX2 mux_inst_1254 (
  .O(mux_o_1254),
  .I0(mux_o_1237),
  .I1(mux_o_1238),
  .S0(dff_q_4)
);
MUX2 mux_inst_1255 (
  .O(mux_o_1255),
  .I0(mux_o_1239),
  .I1(mux_o_1240),
  .S0(dff_q_3)
);
MUX2 mux_inst_1256 (
  .O(mux_o_1256),
  .I0(mux_o_1241),
  .I1(mux_o_1242),
  .S0(dff_q_3)
);
MUX2 mux_inst_1257 (
  .O(mux_o_1257),
  .I0(mux_o_1243),
  .I1(mux_o_1244),
  .S0(dff_q_3)
);
MUX2 mux_inst_1258 (
  .O(mux_o_1258),
  .I0(mux_o_1245),
  .I1(mux_o_1246),
  .S0(dff_q_3)
);
MUX2 mux_inst_1259 (
  .O(mux_o_1259),
  .I0(mux_o_1247),
  .I1(mux_o_1248),
  .S0(dff_q_3)
);
MUX2 mux_inst_1260 (
  .O(mux_o_1260),
  .I0(mux_o_1249),
  .I1(mux_o_1250),
  .S0(dff_q_3)
);
MUX2 mux_inst_1261 (
  .O(mux_o_1261),
  .I0(mux_o_1251),
  .I1(mux_o_1252),
  .S0(dff_q_3)
);
MUX2 mux_inst_1262 (
  .O(mux_o_1262),
  .I0(mux_o_1253),
  .I1(mux_o_1254),
  .S0(dff_q_3)
);
MUX2 mux_inst_1263 (
  .O(mux_o_1263),
  .I0(mux_o_1255),
  .I1(mux_o_1256),
  .S0(dff_q_2)
);
MUX2 mux_inst_1264 (
  .O(mux_o_1264),
  .I0(mux_o_1257),
  .I1(mux_o_1258),
  .S0(dff_q_2)
);
MUX2 mux_inst_1265 (
  .O(mux_o_1265),
  .I0(mux_o_1259),
  .I1(mux_o_1260),
  .S0(dff_q_2)
);
MUX2 mux_inst_1266 (
  .O(mux_o_1266),
  .I0(mux_o_1261),
  .I1(mux_o_1262),
  .S0(dff_q_2)
);
MUX2 mux_inst_1267 (
  .O(mux_o_1267),
  .I0(mux_o_1263),
  .I1(mux_o_1264),
  .S0(dff_q_1)
);
MUX2 mux_inst_1268 (
  .O(mux_o_1268),
  .I0(mux_o_1265),
  .I1(mux_o_1266),
  .S0(dff_q_1)
);
MUX2 mux_inst_1269 (
  .O(dout[9]),
  .I0(mux_o_1267),
  .I1(mux_o_1268),
  .S0(dff_q_0)
);
MUX2 mux_inst_1270 (
  .O(mux_o_1270),
  .I0(sdpb_inst_0_dout[10]),
  .I1(sdpb_inst_1_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1271 (
  .O(mux_o_1271),
  .I0(sdpb_inst_2_dout[10]),
  .I1(sdpb_inst_3_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1272 (
  .O(mux_o_1272),
  .I0(sdpb_inst_4_dout[10]),
  .I1(sdpb_inst_5_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1273 (
  .O(mux_o_1273),
  .I0(sdpb_inst_6_dout[10]),
  .I1(sdpb_inst_7_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1274 (
  .O(mux_o_1274),
  .I0(sdpb_inst_8_dout[10]),
  .I1(sdpb_inst_9_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1275 (
  .O(mux_o_1275),
  .I0(sdpb_inst_10_dout[10]),
  .I1(sdpb_inst_11_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1276 (
  .O(mux_o_1276),
  .I0(sdpb_inst_12_dout[10]),
  .I1(sdpb_inst_13_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1277 (
  .O(mux_o_1277),
  .I0(sdpb_inst_14_dout[10]),
  .I1(sdpb_inst_15_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1278 (
  .O(mux_o_1278),
  .I0(sdpb_inst_16_dout[10]),
  .I1(sdpb_inst_17_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1279 (
  .O(mux_o_1279),
  .I0(sdpb_inst_18_dout[10]),
  .I1(sdpb_inst_19_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1280 (
  .O(mux_o_1280),
  .I0(sdpb_inst_20_dout[10]),
  .I1(sdpb_inst_21_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1281 (
  .O(mux_o_1281),
  .I0(sdpb_inst_22_dout[10]),
  .I1(sdpb_inst_23_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1282 (
  .O(mux_o_1282),
  .I0(sdpb_inst_24_dout[10]),
  .I1(sdpb_inst_25_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1283 (
  .O(mux_o_1283),
  .I0(sdpb_inst_26_dout[10]),
  .I1(sdpb_inst_27_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1284 (
  .O(mux_o_1284),
  .I0(sdpb_inst_28_dout[10]),
  .I1(sdpb_inst_29_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1285 (
  .O(mux_o_1285),
  .I0(sdpb_inst_30_dout[10]),
  .I1(sdpb_inst_31_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1286 (
  .O(mux_o_1286),
  .I0(sdpb_inst_32_dout[10]),
  .I1(sdpb_inst_33_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1287 (
  .O(mux_o_1287),
  .I0(sdpb_inst_34_dout[10]),
  .I1(sdpb_inst_35_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1288 (
  .O(mux_o_1288),
  .I0(sdpb_inst_36_dout[10]),
  .I1(sdpb_inst_37_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1289 (
  .O(mux_o_1289),
  .I0(sdpb_inst_38_dout[10]),
  .I1(sdpb_inst_39_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1290 (
  .O(mux_o_1290),
  .I0(sdpb_inst_40_dout[10]),
  .I1(sdpb_inst_41_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1291 (
  .O(mux_o_1291),
  .I0(sdpb_inst_42_dout[10]),
  .I1(sdpb_inst_43_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1292 (
  .O(mux_o_1292),
  .I0(sdpb_inst_44_dout[10]),
  .I1(sdpb_inst_45_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1293 (
  .O(mux_o_1293),
  .I0(sdpb_inst_46_dout[10]),
  .I1(sdpb_inst_47_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1294 (
  .O(mux_o_1294),
  .I0(sdpb_inst_48_dout[10]),
  .I1(sdpb_inst_49_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1295 (
  .O(mux_o_1295),
  .I0(sdpb_inst_50_dout[10]),
  .I1(sdpb_inst_51_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1296 (
  .O(mux_o_1296),
  .I0(sdpb_inst_52_dout[10]),
  .I1(sdpb_inst_53_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1297 (
  .O(mux_o_1297),
  .I0(sdpb_inst_54_dout[10]),
  .I1(sdpb_inst_55_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1298 (
  .O(mux_o_1298),
  .I0(sdpb_inst_56_dout[10]),
  .I1(sdpb_inst_57_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1299 (
  .O(mux_o_1299),
  .I0(sdpb_inst_58_dout[10]),
  .I1(sdpb_inst_59_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1300 (
  .O(mux_o_1300),
  .I0(sdpb_inst_60_dout[10]),
  .I1(sdpb_inst_61_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1301 (
  .O(mux_o_1301),
  .I0(sdpb_inst_62_dout[10]),
  .I1(sdpb_inst_63_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1302 (
  .O(mux_o_1302),
  .I0(sdpb_inst_64_dout[10]),
  .I1(sdpb_inst_65_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1303 (
  .O(mux_o_1303),
  .I0(sdpb_inst_66_dout[10]),
  .I1(sdpb_inst_67_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1304 (
  .O(mux_o_1304),
  .I0(sdpb_inst_68_dout[10]),
  .I1(sdpb_inst_69_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1305 (
  .O(mux_o_1305),
  .I0(sdpb_inst_70_dout[10]),
  .I1(sdpb_inst_71_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1306 (
  .O(mux_o_1306),
  .I0(sdpb_inst_72_dout[10]),
  .I1(sdpb_inst_73_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1307 (
  .O(mux_o_1307),
  .I0(sdpb_inst_74_dout[10]),
  .I1(sdpb_inst_75_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1308 (
  .O(mux_o_1308),
  .I0(sdpb_inst_76_dout[10]),
  .I1(sdpb_inst_77_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1309 (
  .O(mux_o_1309),
  .I0(sdpb_inst_78_dout[10]),
  .I1(sdpb_inst_79_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1310 (
  .O(mux_o_1310),
  .I0(sdpb_inst_80_dout[10]),
  .I1(sdpb_inst_81_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1311 (
  .O(mux_o_1311),
  .I0(sdpb_inst_82_dout[10]),
  .I1(sdpb_inst_83_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1312 (
  .O(mux_o_1312),
  .I0(sdpb_inst_84_dout[10]),
  .I1(sdpb_inst_85_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1313 (
  .O(mux_o_1313),
  .I0(sdpb_inst_86_dout[10]),
  .I1(sdpb_inst_87_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1314 (
  .O(mux_o_1314),
  .I0(sdpb_inst_88_dout[10]),
  .I1(sdpb_inst_89_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1315 (
  .O(mux_o_1315),
  .I0(sdpb_inst_90_dout[10]),
  .I1(sdpb_inst_91_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1316 (
  .O(mux_o_1316),
  .I0(sdpb_inst_92_dout[10]),
  .I1(sdpb_inst_93_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1317 (
  .O(mux_o_1317),
  .I0(sdpb_inst_94_dout[10]),
  .I1(sdpb_inst_95_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1318 (
  .O(mux_o_1318),
  .I0(sdpb_inst_96_dout[10]),
  .I1(sdpb_inst_97_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1319 (
  .O(mux_o_1319),
  .I0(sdpb_inst_98_dout[10]),
  .I1(sdpb_inst_99_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1320 (
  .O(mux_o_1320),
  .I0(sdpb_inst_100_dout[10]),
  .I1(sdpb_inst_101_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1321 (
  .O(mux_o_1321),
  .I0(sdpb_inst_102_dout[10]),
  .I1(sdpb_inst_103_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1322 (
  .O(mux_o_1322),
  .I0(sdpb_inst_104_dout[10]),
  .I1(sdpb_inst_105_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1323 (
  .O(mux_o_1323),
  .I0(sdpb_inst_106_dout[10]),
  .I1(sdpb_inst_107_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1324 (
  .O(mux_o_1324),
  .I0(sdpb_inst_108_dout[10]),
  .I1(sdpb_inst_109_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1325 (
  .O(mux_o_1325),
  .I0(sdpb_inst_110_dout[10]),
  .I1(sdpb_inst_111_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1326 (
  .O(mux_o_1326),
  .I0(sdpb_inst_112_dout[10]),
  .I1(sdpb_inst_113_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1327 (
  .O(mux_o_1327),
  .I0(sdpb_inst_114_dout[10]),
  .I1(sdpb_inst_115_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1328 (
  .O(mux_o_1328),
  .I0(sdpb_inst_116_dout[10]),
  .I1(sdpb_inst_117_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1329 (
  .O(mux_o_1329),
  .I0(sdpb_inst_118_dout[10]),
  .I1(sdpb_inst_119_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1330 (
  .O(mux_o_1330),
  .I0(sdpb_inst_120_dout[10]),
  .I1(sdpb_inst_121_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1331 (
  .O(mux_o_1331),
  .I0(sdpb_inst_122_dout[10]),
  .I1(sdpb_inst_123_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1332 (
  .O(mux_o_1332),
  .I0(sdpb_inst_124_dout[10]),
  .I1(sdpb_inst_125_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1333 (
  .O(mux_o_1333),
  .I0(sdpb_inst_126_dout[10]),
  .I1(sdpb_inst_127_dout[10]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1334 (
  .O(mux_o_1334),
  .I0(mux_o_1270),
  .I1(mux_o_1271),
  .S0(dff_q_5)
);
MUX2 mux_inst_1335 (
  .O(mux_o_1335),
  .I0(mux_o_1272),
  .I1(mux_o_1273),
  .S0(dff_q_5)
);
MUX2 mux_inst_1336 (
  .O(mux_o_1336),
  .I0(mux_o_1274),
  .I1(mux_o_1275),
  .S0(dff_q_5)
);
MUX2 mux_inst_1337 (
  .O(mux_o_1337),
  .I0(mux_o_1276),
  .I1(mux_o_1277),
  .S0(dff_q_5)
);
MUX2 mux_inst_1338 (
  .O(mux_o_1338),
  .I0(mux_o_1278),
  .I1(mux_o_1279),
  .S0(dff_q_5)
);
MUX2 mux_inst_1339 (
  .O(mux_o_1339),
  .I0(mux_o_1280),
  .I1(mux_o_1281),
  .S0(dff_q_5)
);
MUX2 mux_inst_1340 (
  .O(mux_o_1340),
  .I0(mux_o_1282),
  .I1(mux_o_1283),
  .S0(dff_q_5)
);
MUX2 mux_inst_1341 (
  .O(mux_o_1341),
  .I0(mux_o_1284),
  .I1(mux_o_1285),
  .S0(dff_q_5)
);
MUX2 mux_inst_1342 (
  .O(mux_o_1342),
  .I0(mux_o_1286),
  .I1(mux_o_1287),
  .S0(dff_q_5)
);
MUX2 mux_inst_1343 (
  .O(mux_o_1343),
  .I0(mux_o_1288),
  .I1(mux_o_1289),
  .S0(dff_q_5)
);
MUX2 mux_inst_1344 (
  .O(mux_o_1344),
  .I0(mux_o_1290),
  .I1(mux_o_1291),
  .S0(dff_q_5)
);
MUX2 mux_inst_1345 (
  .O(mux_o_1345),
  .I0(mux_o_1292),
  .I1(mux_o_1293),
  .S0(dff_q_5)
);
MUX2 mux_inst_1346 (
  .O(mux_o_1346),
  .I0(mux_o_1294),
  .I1(mux_o_1295),
  .S0(dff_q_5)
);
MUX2 mux_inst_1347 (
  .O(mux_o_1347),
  .I0(mux_o_1296),
  .I1(mux_o_1297),
  .S0(dff_q_5)
);
MUX2 mux_inst_1348 (
  .O(mux_o_1348),
  .I0(mux_o_1298),
  .I1(mux_o_1299),
  .S0(dff_q_5)
);
MUX2 mux_inst_1349 (
  .O(mux_o_1349),
  .I0(mux_o_1300),
  .I1(mux_o_1301),
  .S0(dff_q_5)
);
MUX2 mux_inst_1350 (
  .O(mux_o_1350),
  .I0(mux_o_1302),
  .I1(mux_o_1303),
  .S0(dff_q_5)
);
MUX2 mux_inst_1351 (
  .O(mux_o_1351),
  .I0(mux_o_1304),
  .I1(mux_o_1305),
  .S0(dff_q_5)
);
MUX2 mux_inst_1352 (
  .O(mux_o_1352),
  .I0(mux_o_1306),
  .I1(mux_o_1307),
  .S0(dff_q_5)
);
MUX2 mux_inst_1353 (
  .O(mux_o_1353),
  .I0(mux_o_1308),
  .I1(mux_o_1309),
  .S0(dff_q_5)
);
MUX2 mux_inst_1354 (
  .O(mux_o_1354),
  .I0(mux_o_1310),
  .I1(mux_o_1311),
  .S0(dff_q_5)
);
MUX2 mux_inst_1355 (
  .O(mux_o_1355),
  .I0(mux_o_1312),
  .I1(mux_o_1313),
  .S0(dff_q_5)
);
MUX2 mux_inst_1356 (
  .O(mux_o_1356),
  .I0(mux_o_1314),
  .I1(mux_o_1315),
  .S0(dff_q_5)
);
MUX2 mux_inst_1357 (
  .O(mux_o_1357),
  .I0(mux_o_1316),
  .I1(mux_o_1317),
  .S0(dff_q_5)
);
MUX2 mux_inst_1358 (
  .O(mux_o_1358),
  .I0(mux_o_1318),
  .I1(mux_o_1319),
  .S0(dff_q_5)
);
MUX2 mux_inst_1359 (
  .O(mux_o_1359),
  .I0(mux_o_1320),
  .I1(mux_o_1321),
  .S0(dff_q_5)
);
MUX2 mux_inst_1360 (
  .O(mux_o_1360),
  .I0(mux_o_1322),
  .I1(mux_o_1323),
  .S0(dff_q_5)
);
MUX2 mux_inst_1361 (
  .O(mux_o_1361),
  .I0(mux_o_1324),
  .I1(mux_o_1325),
  .S0(dff_q_5)
);
MUX2 mux_inst_1362 (
  .O(mux_o_1362),
  .I0(mux_o_1326),
  .I1(mux_o_1327),
  .S0(dff_q_5)
);
MUX2 mux_inst_1363 (
  .O(mux_o_1363),
  .I0(mux_o_1328),
  .I1(mux_o_1329),
  .S0(dff_q_5)
);
MUX2 mux_inst_1364 (
  .O(mux_o_1364),
  .I0(mux_o_1330),
  .I1(mux_o_1331),
  .S0(dff_q_5)
);
MUX2 mux_inst_1365 (
  .O(mux_o_1365),
  .I0(mux_o_1332),
  .I1(mux_o_1333),
  .S0(dff_q_5)
);
MUX2 mux_inst_1366 (
  .O(mux_o_1366),
  .I0(mux_o_1334),
  .I1(mux_o_1335),
  .S0(dff_q_4)
);
MUX2 mux_inst_1367 (
  .O(mux_o_1367),
  .I0(mux_o_1336),
  .I1(mux_o_1337),
  .S0(dff_q_4)
);
MUX2 mux_inst_1368 (
  .O(mux_o_1368),
  .I0(mux_o_1338),
  .I1(mux_o_1339),
  .S0(dff_q_4)
);
MUX2 mux_inst_1369 (
  .O(mux_o_1369),
  .I0(mux_o_1340),
  .I1(mux_o_1341),
  .S0(dff_q_4)
);
MUX2 mux_inst_1370 (
  .O(mux_o_1370),
  .I0(mux_o_1342),
  .I1(mux_o_1343),
  .S0(dff_q_4)
);
MUX2 mux_inst_1371 (
  .O(mux_o_1371),
  .I0(mux_o_1344),
  .I1(mux_o_1345),
  .S0(dff_q_4)
);
MUX2 mux_inst_1372 (
  .O(mux_o_1372),
  .I0(mux_o_1346),
  .I1(mux_o_1347),
  .S0(dff_q_4)
);
MUX2 mux_inst_1373 (
  .O(mux_o_1373),
  .I0(mux_o_1348),
  .I1(mux_o_1349),
  .S0(dff_q_4)
);
MUX2 mux_inst_1374 (
  .O(mux_o_1374),
  .I0(mux_o_1350),
  .I1(mux_o_1351),
  .S0(dff_q_4)
);
MUX2 mux_inst_1375 (
  .O(mux_o_1375),
  .I0(mux_o_1352),
  .I1(mux_o_1353),
  .S0(dff_q_4)
);
MUX2 mux_inst_1376 (
  .O(mux_o_1376),
  .I0(mux_o_1354),
  .I1(mux_o_1355),
  .S0(dff_q_4)
);
MUX2 mux_inst_1377 (
  .O(mux_o_1377),
  .I0(mux_o_1356),
  .I1(mux_o_1357),
  .S0(dff_q_4)
);
MUX2 mux_inst_1378 (
  .O(mux_o_1378),
  .I0(mux_o_1358),
  .I1(mux_o_1359),
  .S0(dff_q_4)
);
MUX2 mux_inst_1379 (
  .O(mux_o_1379),
  .I0(mux_o_1360),
  .I1(mux_o_1361),
  .S0(dff_q_4)
);
MUX2 mux_inst_1380 (
  .O(mux_o_1380),
  .I0(mux_o_1362),
  .I1(mux_o_1363),
  .S0(dff_q_4)
);
MUX2 mux_inst_1381 (
  .O(mux_o_1381),
  .I0(mux_o_1364),
  .I1(mux_o_1365),
  .S0(dff_q_4)
);
MUX2 mux_inst_1382 (
  .O(mux_o_1382),
  .I0(mux_o_1366),
  .I1(mux_o_1367),
  .S0(dff_q_3)
);
MUX2 mux_inst_1383 (
  .O(mux_o_1383),
  .I0(mux_o_1368),
  .I1(mux_o_1369),
  .S0(dff_q_3)
);
MUX2 mux_inst_1384 (
  .O(mux_o_1384),
  .I0(mux_o_1370),
  .I1(mux_o_1371),
  .S0(dff_q_3)
);
MUX2 mux_inst_1385 (
  .O(mux_o_1385),
  .I0(mux_o_1372),
  .I1(mux_o_1373),
  .S0(dff_q_3)
);
MUX2 mux_inst_1386 (
  .O(mux_o_1386),
  .I0(mux_o_1374),
  .I1(mux_o_1375),
  .S0(dff_q_3)
);
MUX2 mux_inst_1387 (
  .O(mux_o_1387),
  .I0(mux_o_1376),
  .I1(mux_o_1377),
  .S0(dff_q_3)
);
MUX2 mux_inst_1388 (
  .O(mux_o_1388),
  .I0(mux_o_1378),
  .I1(mux_o_1379),
  .S0(dff_q_3)
);
MUX2 mux_inst_1389 (
  .O(mux_o_1389),
  .I0(mux_o_1380),
  .I1(mux_o_1381),
  .S0(dff_q_3)
);
MUX2 mux_inst_1390 (
  .O(mux_o_1390),
  .I0(mux_o_1382),
  .I1(mux_o_1383),
  .S0(dff_q_2)
);
MUX2 mux_inst_1391 (
  .O(mux_o_1391),
  .I0(mux_o_1384),
  .I1(mux_o_1385),
  .S0(dff_q_2)
);
MUX2 mux_inst_1392 (
  .O(mux_o_1392),
  .I0(mux_o_1386),
  .I1(mux_o_1387),
  .S0(dff_q_2)
);
MUX2 mux_inst_1393 (
  .O(mux_o_1393),
  .I0(mux_o_1388),
  .I1(mux_o_1389),
  .S0(dff_q_2)
);
MUX2 mux_inst_1394 (
  .O(mux_o_1394),
  .I0(mux_o_1390),
  .I1(mux_o_1391),
  .S0(dff_q_1)
);
MUX2 mux_inst_1395 (
  .O(mux_o_1395),
  .I0(mux_o_1392),
  .I1(mux_o_1393),
  .S0(dff_q_1)
);
MUX2 mux_inst_1396 (
  .O(dout[10]),
  .I0(mux_o_1394),
  .I1(mux_o_1395),
  .S0(dff_q_0)
);
MUX2 mux_inst_1397 (
  .O(mux_o_1397),
  .I0(sdpb_inst_0_dout[11]),
  .I1(sdpb_inst_1_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1398 (
  .O(mux_o_1398),
  .I0(sdpb_inst_2_dout[11]),
  .I1(sdpb_inst_3_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1399 (
  .O(mux_o_1399),
  .I0(sdpb_inst_4_dout[11]),
  .I1(sdpb_inst_5_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1400 (
  .O(mux_o_1400),
  .I0(sdpb_inst_6_dout[11]),
  .I1(sdpb_inst_7_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1401 (
  .O(mux_o_1401),
  .I0(sdpb_inst_8_dout[11]),
  .I1(sdpb_inst_9_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1402 (
  .O(mux_o_1402),
  .I0(sdpb_inst_10_dout[11]),
  .I1(sdpb_inst_11_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1403 (
  .O(mux_o_1403),
  .I0(sdpb_inst_12_dout[11]),
  .I1(sdpb_inst_13_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1404 (
  .O(mux_o_1404),
  .I0(sdpb_inst_14_dout[11]),
  .I1(sdpb_inst_15_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1405 (
  .O(mux_o_1405),
  .I0(sdpb_inst_16_dout[11]),
  .I1(sdpb_inst_17_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1406 (
  .O(mux_o_1406),
  .I0(sdpb_inst_18_dout[11]),
  .I1(sdpb_inst_19_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1407 (
  .O(mux_o_1407),
  .I0(sdpb_inst_20_dout[11]),
  .I1(sdpb_inst_21_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1408 (
  .O(mux_o_1408),
  .I0(sdpb_inst_22_dout[11]),
  .I1(sdpb_inst_23_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1409 (
  .O(mux_o_1409),
  .I0(sdpb_inst_24_dout[11]),
  .I1(sdpb_inst_25_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1410 (
  .O(mux_o_1410),
  .I0(sdpb_inst_26_dout[11]),
  .I1(sdpb_inst_27_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1411 (
  .O(mux_o_1411),
  .I0(sdpb_inst_28_dout[11]),
  .I1(sdpb_inst_29_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1412 (
  .O(mux_o_1412),
  .I0(sdpb_inst_30_dout[11]),
  .I1(sdpb_inst_31_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1413 (
  .O(mux_o_1413),
  .I0(sdpb_inst_32_dout[11]),
  .I1(sdpb_inst_33_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1414 (
  .O(mux_o_1414),
  .I0(sdpb_inst_34_dout[11]),
  .I1(sdpb_inst_35_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1415 (
  .O(mux_o_1415),
  .I0(sdpb_inst_36_dout[11]),
  .I1(sdpb_inst_37_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1416 (
  .O(mux_o_1416),
  .I0(sdpb_inst_38_dout[11]),
  .I1(sdpb_inst_39_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1417 (
  .O(mux_o_1417),
  .I0(sdpb_inst_40_dout[11]),
  .I1(sdpb_inst_41_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1418 (
  .O(mux_o_1418),
  .I0(sdpb_inst_42_dout[11]),
  .I1(sdpb_inst_43_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1419 (
  .O(mux_o_1419),
  .I0(sdpb_inst_44_dout[11]),
  .I1(sdpb_inst_45_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1420 (
  .O(mux_o_1420),
  .I0(sdpb_inst_46_dout[11]),
  .I1(sdpb_inst_47_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1421 (
  .O(mux_o_1421),
  .I0(sdpb_inst_48_dout[11]),
  .I1(sdpb_inst_49_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1422 (
  .O(mux_o_1422),
  .I0(sdpb_inst_50_dout[11]),
  .I1(sdpb_inst_51_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1423 (
  .O(mux_o_1423),
  .I0(sdpb_inst_52_dout[11]),
  .I1(sdpb_inst_53_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1424 (
  .O(mux_o_1424),
  .I0(sdpb_inst_54_dout[11]),
  .I1(sdpb_inst_55_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1425 (
  .O(mux_o_1425),
  .I0(sdpb_inst_56_dout[11]),
  .I1(sdpb_inst_57_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1426 (
  .O(mux_o_1426),
  .I0(sdpb_inst_58_dout[11]),
  .I1(sdpb_inst_59_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1427 (
  .O(mux_o_1427),
  .I0(sdpb_inst_60_dout[11]),
  .I1(sdpb_inst_61_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1428 (
  .O(mux_o_1428),
  .I0(sdpb_inst_62_dout[11]),
  .I1(sdpb_inst_63_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1429 (
  .O(mux_o_1429),
  .I0(sdpb_inst_64_dout[11]),
  .I1(sdpb_inst_65_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1430 (
  .O(mux_o_1430),
  .I0(sdpb_inst_66_dout[11]),
  .I1(sdpb_inst_67_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1431 (
  .O(mux_o_1431),
  .I0(sdpb_inst_68_dout[11]),
  .I1(sdpb_inst_69_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1432 (
  .O(mux_o_1432),
  .I0(sdpb_inst_70_dout[11]),
  .I1(sdpb_inst_71_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1433 (
  .O(mux_o_1433),
  .I0(sdpb_inst_72_dout[11]),
  .I1(sdpb_inst_73_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1434 (
  .O(mux_o_1434),
  .I0(sdpb_inst_74_dout[11]),
  .I1(sdpb_inst_75_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1435 (
  .O(mux_o_1435),
  .I0(sdpb_inst_76_dout[11]),
  .I1(sdpb_inst_77_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1436 (
  .O(mux_o_1436),
  .I0(sdpb_inst_78_dout[11]),
  .I1(sdpb_inst_79_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1437 (
  .O(mux_o_1437),
  .I0(sdpb_inst_80_dout[11]),
  .I1(sdpb_inst_81_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1438 (
  .O(mux_o_1438),
  .I0(sdpb_inst_82_dout[11]),
  .I1(sdpb_inst_83_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1439 (
  .O(mux_o_1439),
  .I0(sdpb_inst_84_dout[11]),
  .I1(sdpb_inst_85_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1440 (
  .O(mux_o_1440),
  .I0(sdpb_inst_86_dout[11]),
  .I1(sdpb_inst_87_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1441 (
  .O(mux_o_1441),
  .I0(sdpb_inst_88_dout[11]),
  .I1(sdpb_inst_89_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1442 (
  .O(mux_o_1442),
  .I0(sdpb_inst_90_dout[11]),
  .I1(sdpb_inst_91_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1443 (
  .O(mux_o_1443),
  .I0(sdpb_inst_92_dout[11]),
  .I1(sdpb_inst_93_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1444 (
  .O(mux_o_1444),
  .I0(sdpb_inst_94_dout[11]),
  .I1(sdpb_inst_95_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1445 (
  .O(mux_o_1445),
  .I0(sdpb_inst_96_dout[11]),
  .I1(sdpb_inst_97_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1446 (
  .O(mux_o_1446),
  .I0(sdpb_inst_98_dout[11]),
  .I1(sdpb_inst_99_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1447 (
  .O(mux_o_1447),
  .I0(sdpb_inst_100_dout[11]),
  .I1(sdpb_inst_101_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1448 (
  .O(mux_o_1448),
  .I0(sdpb_inst_102_dout[11]),
  .I1(sdpb_inst_103_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1449 (
  .O(mux_o_1449),
  .I0(sdpb_inst_104_dout[11]),
  .I1(sdpb_inst_105_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1450 (
  .O(mux_o_1450),
  .I0(sdpb_inst_106_dout[11]),
  .I1(sdpb_inst_107_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1451 (
  .O(mux_o_1451),
  .I0(sdpb_inst_108_dout[11]),
  .I1(sdpb_inst_109_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1452 (
  .O(mux_o_1452),
  .I0(sdpb_inst_110_dout[11]),
  .I1(sdpb_inst_111_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1453 (
  .O(mux_o_1453),
  .I0(sdpb_inst_112_dout[11]),
  .I1(sdpb_inst_113_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1454 (
  .O(mux_o_1454),
  .I0(sdpb_inst_114_dout[11]),
  .I1(sdpb_inst_115_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1455 (
  .O(mux_o_1455),
  .I0(sdpb_inst_116_dout[11]),
  .I1(sdpb_inst_117_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1456 (
  .O(mux_o_1456),
  .I0(sdpb_inst_118_dout[11]),
  .I1(sdpb_inst_119_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1457 (
  .O(mux_o_1457),
  .I0(sdpb_inst_120_dout[11]),
  .I1(sdpb_inst_121_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1458 (
  .O(mux_o_1458),
  .I0(sdpb_inst_122_dout[11]),
  .I1(sdpb_inst_123_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1459 (
  .O(mux_o_1459),
  .I0(sdpb_inst_124_dout[11]),
  .I1(sdpb_inst_125_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1460 (
  .O(mux_o_1460),
  .I0(sdpb_inst_126_dout[11]),
  .I1(sdpb_inst_127_dout[11]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1461 (
  .O(mux_o_1461),
  .I0(mux_o_1397),
  .I1(mux_o_1398),
  .S0(dff_q_5)
);
MUX2 mux_inst_1462 (
  .O(mux_o_1462),
  .I0(mux_o_1399),
  .I1(mux_o_1400),
  .S0(dff_q_5)
);
MUX2 mux_inst_1463 (
  .O(mux_o_1463),
  .I0(mux_o_1401),
  .I1(mux_o_1402),
  .S0(dff_q_5)
);
MUX2 mux_inst_1464 (
  .O(mux_o_1464),
  .I0(mux_o_1403),
  .I1(mux_o_1404),
  .S0(dff_q_5)
);
MUX2 mux_inst_1465 (
  .O(mux_o_1465),
  .I0(mux_o_1405),
  .I1(mux_o_1406),
  .S0(dff_q_5)
);
MUX2 mux_inst_1466 (
  .O(mux_o_1466),
  .I0(mux_o_1407),
  .I1(mux_o_1408),
  .S0(dff_q_5)
);
MUX2 mux_inst_1467 (
  .O(mux_o_1467),
  .I0(mux_o_1409),
  .I1(mux_o_1410),
  .S0(dff_q_5)
);
MUX2 mux_inst_1468 (
  .O(mux_o_1468),
  .I0(mux_o_1411),
  .I1(mux_o_1412),
  .S0(dff_q_5)
);
MUX2 mux_inst_1469 (
  .O(mux_o_1469),
  .I0(mux_o_1413),
  .I1(mux_o_1414),
  .S0(dff_q_5)
);
MUX2 mux_inst_1470 (
  .O(mux_o_1470),
  .I0(mux_o_1415),
  .I1(mux_o_1416),
  .S0(dff_q_5)
);
MUX2 mux_inst_1471 (
  .O(mux_o_1471),
  .I0(mux_o_1417),
  .I1(mux_o_1418),
  .S0(dff_q_5)
);
MUX2 mux_inst_1472 (
  .O(mux_o_1472),
  .I0(mux_o_1419),
  .I1(mux_o_1420),
  .S0(dff_q_5)
);
MUX2 mux_inst_1473 (
  .O(mux_o_1473),
  .I0(mux_o_1421),
  .I1(mux_o_1422),
  .S0(dff_q_5)
);
MUX2 mux_inst_1474 (
  .O(mux_o_1474),
  .I0(mux_o_1423),
  .I1(mux_o_1424),
  .S0(dff_q_5)
);
MUX2 mux_inst_1475 (
  .O(mux_o_1475),
  .I0(mux_o_1425),
  .I1(mux_o_1426),
  .S0(dff_q_5)
);
MUX2 mux_inst_1476 (
  .O(mux_o_1476),
  .I0(mux_o_1427),
  .I1(mux_o_1428),
  .S0(dff_q_5)
);
MUX2 mux_inst_1477 (
  .O(mux_o_1477),
  .I0(mux_o_1429),
  .I1(mux_o_1430),
  .S0(dff_q_5)
);
MUX2 mux_inst_1478 (
  .O(mux_o_1478),
  .I0(mux_o_1431),
  .I1(mux_o_1432),
  .S0(dff_q_5)
);
MUX2 mux_inst_1479 (
  .O(mux_o_1479),
  .I0(mux_o_1433),
  .I1(mux_o_1434),
  .S0(dff_q_5)
);
MUX2 mux_inst_1480 (
  .O(mux_o_1480),
  .I0(mux_o_1435),
  .I1(mux_o_1436),
  .S0(dff_q_5)
);
MUX2 mux_inst_1481 (
  .O(mux_o_1481),
  .I0(mux_o_1437),
  .I1(mux_o_1438),
  .S0(dff_q_5)
);
MUX2 mux_inst_1482 (
  .O(mux_o_1482),
  .I0(mux_o_1439),
  .I1(mux_o_1440),
  .S0(dff_q_5)
);
MUX2 mux_inst_1483 (
  .O(mux_o_1483),
  .I0(mux_o_1441),
  .I1(mux_o_1442),
  .S0(dff_q_5)
);
MUX2 mux_inst_1484 (
  .O(mux_o_1484),
  .I0(mux_o_1443),
  .I1(mux_o_1444),
  .S0(dff_q_5)
);
MUX2 mux_inst_1485 (
  .O(mux_o_1485),
  .I0(mux_o_1445),
  .I1(mux_o_1446),
  .S0(dff_q_5)
);
MUX2 mux_inst_1486 (
  .O(mux_o_1486),
  .I0(mux_o_1447),
  .I1(mux_o_1448),
  .S0(dff_q_5)
);
MUX2 mux_inst_1487 (
  .O(mux_o_1487),
  .I0(mux_o_1449),
  .I1(mux_o_1450),
  .S0(dff_q_5)
);
MUX2 mux_inst_1488 (
  .O(mux_o_1488),
  .I0(mux_o_1451),
  .I1(mux_o_1452),
  .S0(dff_q_5)
);
MUX2 mux_inst_1489 (
  .O(mux_o_1489),
  .I0(mux_o_1453),
  .I1(mux_o_1454),
  .S0(dff_q_5)
);
MUX2 mux_inst_1490 (
  .O(mux_o_1490),
  .I0(mux_o_1455),
  .I1(mux_o_1456),
  .S0(dff_q_5)
);
MUX2 mux_inst_1491 (
  .O(mux_o_1491),
  .I0(mux_o_1457),
  .I1(mux_o_1458),
  .S0(dff_q_5)
);
MUX2 mux_inst_1492 (
  .O(mux_o_1492),
  .I0(mux_o_1459),
  .I1(mux_o_1460),
  .S0(dff_q_5)
);
MUX2 mux_inst_1493 (
  .O(mux_o_1493),
  .I0(mux_o_1461),
  .I1(mux_o_1462),
  .S0(dff_q_4)
);
MUX2 mux_inst_1494 (
  .O(mux_o_1494),
  .I0(mux_o_1463),
  .I1(mux_o_1464),
  .S0(dff_q_4)
);
MUX2 mux_inst_1495 (
  .O(mux_o_1495),
  .I0(mux_o_1465),
  .I1(mux_o_1466),
  .S0(dff_q_4)
);
MUX2 mux_inst_1496 (
  .O(mux_o_1496),
  .I0(mux_o_1467),
  .I1(mux_o_1468),
  .S0(dff_q_4)
);
MUX2 mux_inst_1497 (
  .O(mux_o_1497),
  .I0(mux_o_1469),
  .I1(mux_o_1470),
  .S0(dff_q_4)
);
MUX2 mux_inst_1498 (
  .O(mux_o_1498),
  .I0(mux_o_1471),
  .I1(mux_o_1472),
  .S0(dff_q_4)
);
MUX2 mux_inst_1499 (
  .O(mux_o_1499),
  .I0(mux_o_1473),
  .I1(mux_o_1474),
  .S0(dff_q_4)
);
MUX2 mux_inst_1500 (
  .O(mux_o_1500),
  .I0(mux_o_1475),
  .I1(mux_o_1476),
  .S0(dff_q_4)
);
MUX2 mux_inst_1501 (
  .O(mux_o_1501),
  .I0(mux_o_1477),
  .I1(mux_o_1478),
  .S0(dff_q_4)
);
MUX2 mux_inst_1502 (
  .O(mux_o_1502),
  .I0(mux_o_1479),
  .I1(mux_o_1480),
  .S0(dff_q_4)
);
MUX2 mux_inst_1503 (
  .O(mux_o_1503),
  .I0(mux_o_1481),
  .I1(mux_o_1482),
  .S0(dff_q_4)
);
MUX2 mux_inst_1504 (
  .O(mux_o_1504),
  .I0(mux_o_1483),
  .I1(mux_o_1484),
  .S0(dff_q_4)
);
MUX2 mux_inst_1505 (
  .O(mux_o_1505),
  .I0(mux_o_1485),
  .I1(mux_o_1486),
  .S0(dff_q_4)
);
MUX2 mux_inst_1506 (
  .O(mux_o_1506),
  .I0(mux_o_1487),
  .I1(mux_o_1488),
  .S0(dff_q_4)
);
MUX2 mux_inst_1507 (
  .O(mux_o_1507),
  .I0(mux_o_1489),
  .I1(mux_o_1490),
  .S0(dff_q_4)
);
MUX2 mux_inst_1508 (
  .O(mux_o_1508),
  .I0(mux_o_1491),
  .I1(mux_o_1492),
  .S0(dff_q_4)
);
MUX2 mux_inst_1509 (
  .O(mux_o_1509),
  .I0(mux_o_1493),
  .I1(mux_o_1494),
  .S0(dff_q_3)
);
MUX2 mux_inst_1510 (
  .O(mux_o_1510),
  .I0(mux_o_1495),
  .I1(mux_o_1496),
  .S0(dff_q_3)
);
MUX2 mux_inst_1511 (
  .O(mux_o_1511),
  .I0(mux_o_1497),
  .I1(mux_o_1498),
  .S0(dff_q_3)
);
MUX2 mux_inst_1512 (
  .O(mux_o_1512),
  .I0(mux_o_1499),
  .I1(mux_o_1500),
  .S0(dff_q_3)
);
MUX2 mux_inst_1513 (
  .O(mux_o_1513),
  .I0(mux_o_1501),
  .I1(mux_o_1502),
  .S0(dff_q_3)
);
MUX2 mux_inst_1514 (
  .O(mux_o_1514),
  .I0(mux_o_1503),
  .I1(mux_o_1504),
  .S0(dff_q_3)
);
MUX2 mux_inst_1515 (
  .O(mux_o_1515),
  .I0(mux_o_1505),
  .I1(mux_o_1506),
  .S0(dff_q_3)
);
MUX2 mux_inst_1516 (
  .O(mux_o_1516),
  .I0(mux_o_1507),
  .I1(mux_o_1508),
  .S0(dff_q_3)
);
MUX2 mux_inst_1517 (
  .O(mux_o_1517),
  .I0(mux_o_1509),
  .I1(mux_o_1510),
  .S0(dff_q_2)
);
MUX2 mux_inst_1518 (
  .O(mux_o_1518),
  .I0(mux_o_1511),
  .I1(mux_o_1512),
  .S0(dff_q_2)
);
MUX2 mux_inst_1519 (
  .O(mux_o_1519),
  .I0(mux_o_1513),
  .I1(mux_o_1514),
  .S0(dff_q_2)
);
MUX2 mux_inst_1520 (
  .O(mux_o_1520),
  .I0(mux_o_1515),
  .I1(mux_o_1516),
  .S0(dff_q_2)
);
MUX2 mux_inst_1521 (
  .O(mux_o_1521),
  .I0(mux_o_1517),
  .I1(mux_o_1518),
  .S0(dff_q_1)
);
MUX2 mux_inst_1522 (
  .O(mux_o_1522),
  .I0(mux_o_1519),
  .I1(mux_o_1520),
  .S0(dff_q_1)
);
MUX2 mux_inst_1523 (
  .O(dout[11]),
  .I0(mux_o_1521),
  .I1(mux_o_1522),
  .S0(dff_q_0)
);
MUX2 mux_inst_1524 (
  .O(mux_o_1524),
  .I0(sdpb_inst_0_dout[12]),
  .I1(sdpb_inst_1_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1525 (
  .O(mux_o_1525),
  .I0(sdpb_inst_2_dout[12]),
  .I1(sdpb_inst_3_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1526 (
  .O(mux_o_1526),
  .I0(sdpb_inst_4_dout[12]),
  .I1(sdpb_inst_5_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1527 (
  .O(mux_o_1527),
  .I0(sdpb_inst_6_dout[12]),
  .I1(sdpb_inst_7_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1528 (
  .O(mux_o_1528),
  .I0(sdpb_inst_8_dout[12]),
  .I1(sdpb_inst_9_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1529 (
  .O(mux_o_1529),
  .I0(sdpb_inst_10_dout[12]),
  .I1(sdpb_inst_11_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1530 (
  .O(mux_o_1530),
  .I0(sdpb_inst_12_dout[12]),
  .I1(sdpb_inst_13_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1531 (
  .O(mux_o_1531),
  .I0(sdpb_inst_14_dout[12]),
  .I1(sdpb_inst_15_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1532 (
  .O(mux_o_1532),
  .I0(sdpb_inst_16_dout[12]),
  .I1(sdpb_inst_17_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1533 (
  .O(mux_o_1533),
  .I0(sdpb_inst_18_dout[12]),
  .I1(sdpb_inst_19_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1534 (
  .O(mux_o_1534),
  .I0(sdpb_inst_20_dout[12]),
  .I1(sdpb_inst_21_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1535 (
  .O(mux_o_1535),
  .I0(sdpb_inst_22_dout[12]),
  .I1(sdpb_inst_23_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1536 (
  .O(mux_o_1536),
  .I0(sdpb_inst_24_dout[12]),
  .I1(sdpb_inst_25_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1537 (
  .O(mux_o_1537),
  .I0(sdpb_inst_26_dout[12]),
  .I1(sdpb_inst_27_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1538 (
  .O(mux_o_1538),
  .I0(sdpb_inst_28_dout[12]),
  .I1(sdpb_inst_29_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1539 (
  .O(mux_o_1539),
  .I0(sdpb_inst_30_dout[12]),
  .I1(sdpb_inst_31_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1540 (
  .O(mux_o_1540),
  .I0(sdpb_inst_32_dout[12]),
  .I1(sdpb_inst_33_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1541 (
  .O(mux_o_1541),
  .I0(sdpb_inst_34_dout[12]),
  .I1(sdpb_inst_35_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1542 (
  .O(mux_o_1542),
  .I0(sdpb_inst_36_dout[12]),
  .I1(sdpb_inst_37_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1543 (
  .O(mux_o_1543),
  .I0(sdpb_inst_38_dout[12]),
  .I1(sdpb_inst_39_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1544 (
  .O(mux_o_1544),
  .I0(sdpb_inst_40_dout[12]),
  .I1(sdpb_inst_41_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1545 (
  .O(mux_o_1545),
  .I0(sdpb_inst_42_dout[12]),
  .I1(sdpb_inst_43_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1546 (
  .O(mux_o_1546),
  .I0(sdpb_inst_44_dout[12]),
  .I1(sdpb_inst_45_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1547 (
  .O(mux_o_1547),
  .I0(sdpb_inst_46_dout[12]),
  .I1(sdpb_inst_47_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1548 (
  .O(mux_o_1548),
  .I0(sdpb_inst_48_dout[12]),
  .I1(sdpb_inst_49_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1549 (
  .O(mux_o_1549),
  .I0(sdpb_inst_50_dout[12]),
  .I1(sdpb_inst_51_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1550 (
  .O(mux_o_1550),
  .I0(sdpb_inst_52_dout[12]),
  .I1(sdpb_inst_53_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1551 (
  .O(mux_o_1551),
  .I0(sdpb_inst_54_dout[12]),
  .I1(sdpb_inst_55_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1552 (
  .O(mux_o_1552),
  .I0(sdpb_inst_56_dout[12]),
  .I1(sdpb_inst_57_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1553 (
  .O(mux_o_1553),
  .I0(sdpb_inst_58_dout[12]),
  .I1(sdpb_inst_59_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1554 (
  .O(mux_o_1554),
  .I0(sdpb_inst_60_dout[12]),
  .I1(sdpb_inst_61_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1555 (
  .O(mux_o_1555),
  .I0(sdpb_inst_62_dout[12]),
  .I1(sdpb_inst_63_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1556 (
  .O(mux_o_1556),
  .I0(sdpb_inst_64_dout[12]),
  .I1(sdpb_inst_65_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1557 (
  .O(mux_o_1557),
  .I0(sdpb_inst_66_dout[12]),
  .I1(sdpb_inst_67_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1558 (
  .O(mux_o_1558),
  .I0(sdpb_inst_68_dout[12]),
  .I1(sdpb_inst_69_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1559 (
  .O(mux_o_1559),
  .I0(sdpb_inst_70_dout[12]),
  .I1(sdpb_inst_71_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1560 (
  .O(mux_o_1560),
  .I0(sdpb_inst_72_dout[12]),
  .I1(sdpb_inst_73_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1561 (
  .O(mux_o_1561),
  .I0(sdpb_inst_74_dout[12]),
  .I1(sdpb_inst_75_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1562 (
  .O(mux_o_1562),
  .I0(sdpb_inst_76_dout[12]),
  .I1(sdpb_inst_77_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1563 (
  .O(mux_o_1563),
  .I0(sdpb_inst_78_dout[12]),
  .I1(sdpb_inst_79_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1564 (
  .O(mux_o_1564),
  .I0(sdpb_inst_80_dout[12]),
  .I1(sdpb_inst_81_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1565 (
  .O(mux_o_1565),
  .I0(sdpb_inst_82_dout[12]),
  .I1(sdpb_inst_83_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1566 (
  .O(mux_o_1566),
  .I0(sdpb_inst_84_dout[12]),
  .I1(sdpb_inst_85_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1567 (
  .O(mux_o_1567),
  .I0(sdpb_inst_86_dout[12]),
  .I1(sdpb_inst_87_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1568 (
  .O(mux_o_1568),
  .I0(sdpb_inst_88_dout[12]),
  .I1(sdpb_inst_89_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1569 (
  .O(mux_o_1569),
  .I0(sdpb_inst_90_dout[12]),
  .I1(sdpb_inst_91_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1570 (
  .O(mux_o_1570),
  .I0(sdpb_inst_92_dout[12]),
  .I1(sdpb_inst_93_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1571 (
  .O(mux_o_1571),
  .I0(sdpb_inst_94_dout[12]),
  .I1(sdpb_inst_95_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1572 (
  .O(mux_o_1572),
  .I0(sdpb_inst_96_dout[12]),
  .I1(sdpb_inst_97_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1573 (
  .O(mux_o_1573),
  .I0(sdpb_inst_98_dout[12]),
  .I1(sdpb_inst_99_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1574 (
  .O(mux_o_1574),
  .I0(sdpb_inst_100_dout[12]),
  .I1(sdpb_inst_101_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1575 (
  .O(mux_o_1575),
  .I0(sdpb_inst_102_dout[12]),
  .I1(sdpb_inst_103_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1576 (
  .O(mux_o_1576),
  .I0(sdpb_inst_104_dout[12]),
  .I1(sdpb_inst_105_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1577 (
  .O(mux_o_1577),
  .I0(sdpb_inst_106_dout[12]),
  .I1(sdpb_inst_107_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1578 (
  .O(mux_o_1578),
  .I0(sdpb_inst_108_dout[12]),
  .I1(sdpb_inst_109_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1579 (
  .O(mux_o_1579),
  .I0(sdpb_inst_110_dout[12]),
  .I1(sdpb_inst_111_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1580 (
  .O(mux_o_1580),
  .I0(sdpb_inst_112_dout[12]),
  .I1(sdpb_inst_113_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1581 (
  .O(mux_o_1581),
  .I0(sdpb_inst_114_dout[12]),
  .I1(sdpb_inst_115_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1582 (
  .O(mux_o_1582),
  .I0(sdpb_inst_116_dout[12]),
  .I1(sdpb_inst_117_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1583 (
  .O(mux_o_1583),
  .I0(sdpb_inst_118_dout[12]),
  .I1(sdpb_inst_119_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1584 (
  .O(mux_o_1584),
  .I0(sdpb_inst_120_dout[12]),
  .I1(sdpb_inst_121_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1585 (
  .O(mux_o_1585),
  .I0(sdpb_inst_122_dout[12]),
  .I1(sdpb_inst_123_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1586 (
  .O(mux_o_1586),
  .I0(sdpb_inst_124_dout[12]),
  .I1(sdpb_inst_125_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1587 (
  .O(mux_o_1587),
  .I0(sdpb_inst_126_dout[12]),
  .I1(sdpb_inst_127_dout[12]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1588 (
  .O(mux_o_1588),
  .I0(mux_o_1524),
  .I1(mux_o_1525),
  .S0(dff_q_5)
);
MUX2 mux_inst_1589 (
  .O(mux_o_1589),
  .I0(mux_o_1526),
  .I1(mux_o_1527),
  .S0(dff_q_5)
);
MUX2 mux_inst_1590 (
  .O(mux_o_1590),
  .I0(mux_o_1528),
  .I1(mux_o_1529),
  .S0(dff_q_5)
);
MUX2 mux_inst_1591 (
  .O(mux_o_1591),
  .I0(mux_o_1530),
  .I1(mux_o_1531),
  .S0(dff_q_5)
);
MUX2 mux_inst_1592 (
  .O(mux_o_1592),
  .I0(mux_o_1532),
  .I1(mux_o_1533),
  .S0(dff_q_5)
);
MUX2 mux_inst_1593 (
  .O(mux_o_1593),
  .I0(mux_o_1534),
  .I1(mux_o_1535),
  .S0(dff_q_5)
);
MUX2 mux_inst_1594 (
  .O(mux_o_1594),
  .I0(mux_o_1536),
  .I1(mux_o_1537),
  .S0(dff_q_5)
);
MUX2 mux_inst_1595 (
  .O(mux_o_1595),
  .I0(mux_o_1538),
  .I1(mux_o_1539),
  .S0(dff_q_5)
);
MUX2 mux_inst_1596 (
  .O(mux_o_1596),
  .I0(mux_o_1540),
  .I1(mux_o_1541),
  .S0(dff_q_5)
);
MUX2 mux_inst_1597 (
  .O(mux_o_1597),
  .I0(mux_o_1542),
  .I1(mux_o_1543),
  .S0(dff_q_5)
);
MUX2 mux_inst_1598 (
  .O(mux_o_1598),
  .I0(mux_o_1544),
  .I1(mux_o_1545),
  .S0(dff_q_5)
);
MUX2 mux_inst_1599 (
  .O(mux_o_1599),
  .I0(mux_o_1546),
  .I1(mux_o_1547),
  .S0(dff_q_5)
);
MUX2 mux_inst_1600 (
  .O(mux_o_1600),
  .I0(mux_o_1548),
  .I1(mux_o_1549),
  .S0(dff_q_5)
);
MUX2 mux_inst_1601 (
  .O(mux_o_1601),
  .I0(mux_o_1550),
  .I1(mux_o_1551),
  .S0(dff_q_5)
);
MUX2 mux_inst_1602 (
  .O(mux_o_1602),
  .I0(mux_o_1552),
  .I1(mux_o_1553),
  .S0(dff_q_5)
);
MUX2 mux_inst_1603 (
  .O(mux_o_1603),
  .I0(mux_o_1554),
  .I1(mux_o_1555),
  .S0(dff_q_5)
);
MUX2 mux_inst_1604 (
  .O(mux_o_1604),
  .I0(mux_o_1556),
  .I1(mux_o_1557),
  .S0(dff_q_5)
);
MUX2 mux_inst_1605 (
  .O(mux_o_1605),
  .I0(mux_o_1558),
  .I1(mux_o_1559),
  .S0(dff_q_5)
);
MUX2 mux_inst_1606 (
  .O(mux_o_1606),
  .I0(mux_o_1560),
  .I1(mux_o_1561),
  .S0(dff_q_5)
);
MUX2 mux_inst_1607 (
  .O(mux_o_1607),
  .I0(mux_o_1562),
  .I1(mux_o_1563),
  .S0(dff_q_5)
);
MUX2 mux_inst_1608 (
  .O(mux_o_1608),
  .I0(mux_o_1564),
  .I1(mux_o_1565),
  .S0(dff_q_5)
);
MUX2 mux_inst_1609 (
  .O(mux_o_1609),
  .I0(mux_o_1566),
  .I1(mux_o_1567),
  .S0(dff_q_5)
);
MUX2 mux_inst_1610 (
  .O(mux_o_1610),
  .I0(mux_o_1568),
  .I1(mux_o_1569),
  .S0(dff_q_5)
);
MUX2 mux_inst_1611 (
  .O(mux_o_1611),
  .I0(mux_o_1570),
  .I1(mux_o_1571),
  .S0(dff_q_5)
);
MUX2 mux_inst_1612 (
  .O(mux_o_1612),
  .I0(mux_o_1572),
  .I1(mux_o_1573),
  .S0(dff_q_5)
);
MUX2 mux_inst_1613 (
  .O(mux_o_1613),
  .I0(mux_o_1574),
  .I1(mux_o_1575),
  .S0(dff_q_5)
);
MUX2 mux_inst_1614 (
  .O(mux_o_1614),
  .I0(mux_o_1576),
  .I1(mux_o_1577),
  .S0(dff_q_5)
);
MUX2 mux_inst_1615 (
  .O(mux_o_1615),
  .I0(mux_o_1578),
  .I1(mux_o_1579),
  .S0(dff_q_5)
);
MUX2 mux_inst_1616 (
  .O(mux_o_1616),
  .I0(mux_o_1580),
  .I1(mux_o_1581),
  .S0(dff_q_5)
);
MUX2 mux_inst_1617 (
  .O(mux_o_1617),
  .I0(mux_o_1582),
  .I1(mux_o_1583),
  .S0(dff_q_5)
);
MUX2 mux_inst_1618 (
  .O(mux_o_1618),
  .I0(mux_o_1584),
  .I1(mux_o_1585),
  .S0(dff_q_5)
);
MUX2 mux_inst_1619 (
  .O(mux_o_1619),
  .I0(mux_o_1586),
  .I1(mux_o_1587),
  .S0(dff_q_5)
);
MUX2 mux_inst_1620 (
  .O(mux_o_1620),
  .I0(mux_o_1588),
  .I1(mux_o_1589),
  .S0(dff_q_4)
);
MUX2 mux_inst_1621 (
  .O(mux_o_1621),
  .I0(mux_o_1590),
  .I1(mux_o_1591),
  .S0(dff_q_4)
);
MUX2 mux_inst_1622 (
  .O(mux_o_1622),
  .I0(mux_o_1592),
  .I1(mux_o_1593),
  .S0(dff_q_4)
);
MUX2 mux_inst_1623 (
  .O(mux_o_1623),
  .I0(mux_o_1594),
  .I1(mux_o_1595),
  .S0(dff_q_4)
);
MUX2 mux_inst_1624 (
  .O(mux_o_1624),
  .I0(mux_o_1596),
  .I1(mux_o_1597),
  .S0(dff_q_4)
);
MUX2 mux_inst_1625 (
  .O(mux_o_1625),
  .I0(mux_o_1598),
  .I1(mux_o_1599),
  .S0(dff_q_4)
);
MUX2 mux_inst_1626 (
  .O(mux_o_1626),
  .I0(mux_o_1600),
  .I1(mux_o_1601),
  .S0(dff_q_4)
);
MUX2 mux_inst_1627 (
  .O(mux_o_1627),
  .I0(mux_o_1602),
  .I1(mux_o_1603),
  .S0(dff_q_4)
);
MUX2 mux_inst_1628 (
  .O(mux_o_1628),
  .I0(mux_o_1604),
  .I1(mux_o_1605),
  .S0(dff_q_4)
);
MUX2 mux_inst_1629 (
  .O(mux_o_1629),
  .I0(mux_o_1606),
  .I1(mux_o_1607),
  .S0(dff_q_4)
);
MUX2 mux_inst_1630 (
  .O(mux_o_1630),
  .I0(mux_o_1608),
  .I1(mux_o_1609),
  .S0(dff_q_4)
);
MUX2 mux_inst_1631 (
  .O(mux_o_1631),
  .I0(mux_o_1610),
  .I1(mux_o_1611),
  .S0(dff_q_4)
);
MUX2 mux_inst_1632 (
  .O(mux_o_1632),
  .I0(mux_o_1612),
  .I1(mux_o_1613),
  .S0(dff_q_4)
);
MUX2 mux_inst_1633 (
  .O(mux_o_1633),
  .I0(mux_o_1614),
  .I1(mux_o_1615),
  .S0(dff_q_4)
);
MUX2 mux_inst_1634 (
  .O(mux_o_1634),
  .I0(mux_o_1616),
  .I1(mux_o_1617),
  .S0(dff_q_4)
);
MUX2 mux_inst_1635 (
  .O(mux_o_1635),
  .I0(mux_o_1618),
  .I1(mux_o_1619),
  .S0(dff_q_4)
);
MUX2 mux_inst_1636 (
  .O(mux_o_1636),
  .I0(mux_o_1620),
  .I1(mux_o_1621),
  .S0(dff_q_3)
);
MUX2 mux_inst_1637 (
  .O(mux_o_1637),
  .I0(mux_o_1622),
  .I1(mux_o_1623),
  .S0(dff_q_3)
);
MUX2 mux_inst_1638 (
  .O(mux_o_1638),
  .I0(mux_o_1624),
  .I1(mux_o_1625),
  .S0(dff_q_3)
);
MUX2 mux_inst_1639 (
  .O(mux_o_1639),
  .I0(mux_o_1626),
  .I1(mux_o_1627),
  .S0(dff_q_3)
);
MUX2 mux_inst_1640 (
  .O(mux_o_1640),
  .I0(mux_o_1628),
  .I1(mux_o_1629),
  .S0(dff_q_3)
);
MUX2 mux_inst_1641 (
  .O(mux_o_1641),
  .I0(mux_o_1630),
  .I1(mux_o_1631),
  .S0(dff_q_3)
);
MUX2 mux_inst_1642 (
  .O(mux_o_1642),
  .I0(mux_o_1632),
  .I1(mux_o_1633),
  .S0(dff_q_3)
);
MUX2 mux_inst_1643 (
  .O(mux_o_1643),
  .I0(mux_o_1634),
  .I1(mux_o_1635),
  .S0(dff_q_3)
);
MUX2 mux_inst_1644 (
  .O(mux_o_1644),
  .I0(mux_o_1636),
  .I1(mux_o_1637),
  .S0(dff_q_2)
);
MUX2 mux_inst_1645 (
  .O(mux_o_1645),
  .I0(mux_o_1638),
  .I1(mux_o_1639),
  .S0(dff_q_2)
);
MUX2 mux_inst_1646 (
  .O(mux_o_1646),
  .I0(mux_o_1640),
  .I1(mux_o_1641),
  .S0(dff_q_2)
);
MUX2 mux_inst_1647 (
  .O(mux_o_1647),
  .I0(mux_o_1642),
  .I1(mux_o_1643),
  .S0(dff_q_2)
);
MUX2 mux_inst_1648 (
  .O(mux_o_1648),
  .I0(mux_o_1644),
  .I1(mux_o_1645),
  .S0(dff_q_1)
);
MUX2 mux_inst_1649 (
  .O(mux_o_1649),
  .I0(mux_o_1646),
  .I1(mux_o_1647),
  .S0(dff_q_1)
);
MUX2 mux_inst_1650 (
  .O(dout[12]),
  .I0(mux_o_1648),
  .I1(mux_o_1649),
  .S0(dff_q_0)
);
MUX2 mux_inst_1651 (
  .O(mux_o_1651),
  .I0(sdpb_inst_0_dout[13]),
  .I1(sdpb_inst_1_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1652 (
  .O(mux_o_1652),
  .I0(sdpb_inst_2_dout[13]),
  .I1(sdpb_inst_3_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1653 (
  .O(mux_o_1653),
  .I0(sdpb_inst_4_dout[13]),
  .I1(sdpb_inst_5_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1654 (
  .O(mux_o_1654),
  .I0(sdpb_inst_6_dout[13]),
  .I1(sdpb_inst_7_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1655 (
  .O(mux_o_1655),
  .I0(sdpb_inst_8_dout[13]),
  .I1(sdpb_inst_9_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1656 (
  .O(mux_o_1656),
  .I0(sdpb_inst_10_dout[13]),
  .I1(sdpb_inst_11_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1657 (
  .O(mux_o_1657),
  .I0(sdpb_inst_12_dout[13]),
  .I1(sdpb_inst_13_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1658 (
  .O(mux_o_1658),
  .I0(sdpb_inst_14_dout[13]),
  .I1(sdpb_inst_15_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1659 (
  .O(mux_o_1659),
  .I0(sdpb_inst_16_dout[13]),
  .I1(sdpb_inst_17_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1660 (
  .O(mux_o_1660),
  .I0(sdpb_inst_18_dout[13]),
  .I1(sdpb_inst_19_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1661 (
  .O(mux_o_1661),
  .I0(sdpb_inst_20_dout[13]),
  .I1(sdpb_inst_21_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1662 (
  .O(mux_o_1662),
  .I0(sdpb_inst_22_dout[13]),
  .I1(sdpb_inst_23_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1663 (
  .O(mux_o_1663),
  .I0(sdpb_inst_24_dout[13]),
  .I1(sdpb_inst_25_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1664 (
  .O(mux_o_1664),
  .I0(sdpb_inst_26_dout[13]),
  .I1(sdpb_inst_27_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1665 (
  .O(mux_o_1665),
  .I0(sdpb_inst_28_dout[13]),
  .I1(sdpb_inst_29_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1666 (
  .O(mux_o_1666),
  .I0(sdpb_inst_30_dout[13]),
  .I1(sdpb_inst_31_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1667 (
  .O(mux_o_1667),
  .I0(sdpb_inst_32_dout[13]),
  .I1(sdpb_inst_33_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1668 (
  .O(mux_o_1668),
  .I0(sdpb_inst_34_dout[13]),
  .I1(sdpb_inst_35_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1669 (
  .O(mux_o_1669),
  .I0(sdpb_inst_36_dout[13]),
  .I1(sdpb_inst_37_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1670 (
  .O(mux_o_1670),
  .I0(sdpb_inst_38_dout[13]),
  .I1(sdpb_inst_39_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1671 (
  .O(mux_o_1671),
  .I0(sdpb_inst_40_dout[13]),
  .I1(sdpb_inst_41_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1672 (
  .O(mux_o_1672),
  .I0(sdpb_inst_42_dout[13]),
  .I1(sdpb_inst_43_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1673 (
  .O(mux_o_1673),
  .I0(sdpb_inst_44_dout[13]),
  .I1(sdpb_inst_45_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1674 (
  .O(mux_o_1674),
  .I0(sdpb_inst_46_dout[13]),
  .I1(sdpb_inst_47_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1675 (
  .O(mux_o_1675),
  .I0(sdpb_inst_48_dout[13]),
  .I1(sdpb_inst_49_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1676 (
  .O(mux_o_1676),
  .I0(sdpb_inst_50_dout[13]),
  .I1(sdpb_inst_51_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1677 (
  .O(mux_o_1677),
  .I0(sdpb_inst_52_dout[13]),
  .I1(sdpb_inst_53_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1678 (
  .O(mux_o_1678),
  .I0(sdpb_inst_54_dout[13]),
  .I1(sdpb_inst_55_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1679 (
  .O(mux_o_1679),
  .I0(sdpb_inst_56_dout[13]),
  .I1(sdpb_inst_57_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1680 (
  .O(mux_o_1680),
  .I0(sdpb_inst_58_dout[13]),
  .I1(sdpb_inst_59_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1681 (
  .O(mux_o_1681),
  .I0(sdpb_inst_60_dout[13]),
  .I1(sdpb_inst_61_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1682 (
  .O(mux_o_1682),
  .I0(sdpb_inst_62_dout[13]),
  .I1(sdpb_inst_63_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1683 (
  .O(mux_o_1683),
  .I0(sdpb_inst_64_dout[13]),
  .I1(sdpb_inst_65_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1684 (
  .O(mux_o_1684),
  .I0(sdpb_inst_66_dout[13]),
  .I1(sdpb_inst_67_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1685 (
  .O(mux_o_1685),
  .I0(sdpb_inst_68_dout[13]),
  .I1(sdpb_inst_69_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1686 (
  .O(mux_o_1686),
  .I0(sdpb_inst_70_dout[13]),
  .I1(sdpb_inst_71_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1687 (
  .O(mux_o_1687),
  .I0(sdpb_inst_72_dout[13]),
  .I1(sdpb_inst_73_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1688 (
  .O(mux_o_1688),
  .I0(sdpb_inst_74_dout[13]),
  .I1(sdpb_inst_75_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1689 (
  .O(mux_o_1689),
  .I0(sdpb_inst_76_dout[13]),
  .I1(sdpb_inst_77_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1690 (
  .O(mux_o_1690),
  .I0(sdpb_inst_78_dout[13]),
  .I1(sdpb_inst_79_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1691 (
  .O(mux_o_1691),
  .I0(sdpb_inst_80_dout[13]),
  .I1(sdpb_inst_81_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1692 (
  .O(mux_o_1692),
  .I0(sdpb_inst_82_dout[13]),
  .I1(sdpb_inst_83_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1693 (
  .O(mux_o_1693),
  .I0(sdpb_inst_84_dout[13]),
  .I1(sdpb_inst_85_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1694 (
  .O(mux_o_1694),
  .I0(sdpb_inst_86_dout[13]),
  .I1(sdpb_inst_87_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1695 (
  .O(mux_o_1695),
  .I0(sdpb_inst_88_dout[13]),
  .I1(sdpb_inst_89_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1696 (
  .O(mux_o_1696),
  .I0(sdpb_inst_90_dout[13]),
  .I1(sdpb_inst_91_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1697 (
  .O(mux_o_1697),
  .I0(sdpb_inst_92_dout[13]),
  .I1(sdpb_inst_93_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1698 (
  .O(mux_o_1698),
  .I0(sdpb_inst_94_dout[13]),
  .I1(sdpb_inst_95_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1699 (
  .O(mux_o_1699),
  .I0(sdpb_inst_96_dout[13]),
  .I1(sdpb_inst_97_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1700 (
  .O(mux_o_1700),
  .I0(sdpb_inst_98_dout[13]),
  .I1(sdpb_inst_99_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1701 (
  .O(mux_o_1701),
  .I0(sdpb_inst_100_dout[13]),
  .I1(sdpb_inst_101_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1702 (
  .O(mux_o_1702),
  .I0(sdpb_inst_102_dout[13]),
  .I1(sdpb_inst_103_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1703 (
  .O(mux_o_1703),
  .I0(sdpb_inst_104_dout[13]),
  .I1(sdpb_inst_105_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1704 (
  .O(mux_o_1704),
  .I0(sdpb_inst_106_dout[13]),
  .I1(sdpb_inst_107_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1705 (
  .O(mux_o_1705),
  .I0(sdpb_inst_108_dout[13]),
  .I1(sdpb_inst_109_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1706 (
  .O(mux_o_1706),
  .I0(sdpb_inst_110_dout[13]),
  .I1(sdpb_inst_111_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1707 (
  .O(mux_o_1707),
  .I0(sdpb_inst_112_dout[13]),
  .I1(sdpb_inst_113_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1708 (
  .O(mux_o_1708),
  .I0(sdpb_inst_114_dout[13]),
  .I1(sdpb_inst_115_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1709 (
  .O(mux_o_1709),
  .I0(sdpb_inst_116_dout[13]),
  .I1(sdpb_inst_117_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1710 (
  .O(mux_o_1710),
  .I0(sdpb_inst_118_dout[13]),
  .I1(sdpb_inst_119_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1711 (
  .O(mux_o_1711),
  .I0(sdpb_inst_120_dout[13]),
  .I1(sdpb_inst_121_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1712 (
  .O(mux_o_1712),
  .I0(sdpb_inst_122_dout[13]),
  .I1(sdpb_inst_123_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1713 (
  .O(mux_o_1713),
  .I0(sdpb_inst_124_dout[13]),
  .I1(sdpb_inst_125_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1714 (
  .O(mux_o_1714),
  .I0(sdpb_inst_126_dout[13]),
  .I1(sdpb_inst_127_dout[13]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1715 (
  .O(mux_o_1715),
  .I0(mux_o_1651),
  .I1(mux_o_1652),
  .S0(dff_q_5)
);
MUX2 mux_inst_1716 (
  .O(mux_o_1716),
  .I0(mux_o_1653),
  .I1(mux_o_1654),
  .S0(dff_q_5)
);
MUX2 mux_inst_1717 (
  .O(mux_o_1717),
  .I0(mux_o_1655),
  .I1(mux_o_1656),
  .S0(dff_q_5)
);
MUX2 mux_inst_1718 (
  .O(mux_o_1718),
  .I0(mux_o_1657),
  .I1(mux_o_1658),
  .S0(dff_q_5)
);
MUX2 mux_inst_1719 (
  .O(mux_o_1719),
  .I0(mux_o_1659),
  .I1(mux_o_1660),
  .S0(dff_q_5)
);
MUX2 mux_inst_1720 (
  .O(mux_o_1720),
  .I0(mux_o_1661),
  .I1(mux_o_1662),
  .S0(dff_q_5)
);
MUX2 mux_inst_1721 (
  .O(mux_o_1721),
  .I0(mux_o_1663),
  .I1(mux_o_1664),
  .S0(dff_q_5)
);
MUX2 mux_inst_1722 (
  .O(mux_o_1722),
  .I0(mux_o_1665),
  .I1(mux_o_1666),
  .S0(dff_q_5)
);
MUX2 mux_inst_1723 (
  .O(mux_o_1723),
  .I0(mux_o_1667),
  .I1(mux_o_1668),
  .S0(dff_q_5)
);
MUX2 mux_inst_1724 (
  .O(mux_o_1724),
  .I0(mux_o_1669),
  .I1(mux_o_1670),
  .S0(dff_q_5)
);
MUX2 mux_inst_1725 (
  .O(mux_o_1725),
  .I0(mux_o_1671),
  .I1(mux_o_1672),
  .S0(dff_q_5)
);
MUX2 mux_inst_1726 (
  .O(mux_o_1726),
  .I0(mux_o_1673),
  .I1(mux_o_1674),
  .S0(dff_q_5)
);
MUX2 mux_inst_1727 (
  .O(mux_o_1727),
  .I0(mux_o_1675),
  .I1(mux_o_1676),
  .S0(dff_q_5)
);
MUX2 mux_inst_1728 (
  .O(mux_o_1728),
  .I0(mux_o_1677),
  .I1(mux_o_1678),
  .S0(dff_q_5)
);
MUX2 mux_inst_1729 (
  .O(mux_o_1729),
  .I0(mux_o_1679),
  .I1(mux_o_1680),
  .S0(dff_q_5)
);
MUX2 mux_inst_1730 (
  .O(mux_o_1730),
  .I0(mux_o_1681),
  .I1(mux_o_1682),
  .S0(dff_q_5)
);
MUX2 mux_inst_1731 (
  .O(mux_o_1731),
  .I0(mux_o_1683),
  .I1(mux_o_1684),
  .S0(dff_q_5)
);
MUX2 mux_inst_1732 (
  .O(mux_o_1732),
  .I0(mux_o_1685),
  .I1(mux_o_1686),
  .S0(dff_q_5)
);
MUX2 mux_inst_1733 (
  .O(mux_o_1733),
  .I0(mux_o_1687),
  .I1(mux_o_1688),
  .S0(dff_q_5)
);
MUX2 mux_inst_1734 (
  .O(mux_o_1734),
  .I0(mux_o_1689),
  .I1(mux_o_1690),
  .S0(dff_q_5)
);
MUX2 mux_inst_1735 (
  .O(mux_o_1735),
  .I0(mux_o_1691),
  .I1(mux_o_1692),
  .S0(dff_q_5)
);
MUX2 mux_inst_1736 (
  .O(mux_o_1736),
  .I0(mux_o_1693),
  .I1(mux_o_1694),
  .S0(dff_q_5)
);
MUX2 mux_inst_1737 (
  .O(mux_o_1737),
  .I0(mux_o_1695),
  .I1(mux_o_1696),
  .S0(dff_q_5)
);
MUX2 mux_inst_1738 (
  .O(mux_o_1738),
  .I0(mux_o_1697),
  .I1(mux_o_1698),
  .S0(dff_q_5)
);
MUX2 mux_inst_1739 (
  .O(mux_o_1739),
  .I0(mux_o_1699),
  .I1(mux_o_1700),
  .S0(dff_q_5)
);
MUX2 mux_inst_1740 (
  .O(mux_o_1740),
  .I0(mux_o_1701),
  .I1(mux_o_1702),
  .S0(dff_q_5)
);
MUX2 mux_inst_1741 (
  .O(mux_o_1741),
  .I0(mux_o_1703),
  .I1(mux_o_1704),
  .S0(dff_q_5)
);
MUX2 mux_inst_1742 (
  .O(mux_o_1742),
  .I0(mux_o_1705),
  .I1(mux_o_1706),
  .S0(dff_q_5)
);
MUX2 mux_inst_1743 (
  .O(mux_o_1743),
  .I0(mux_o_1707),
  .I1(mux_o_1708),
  .S0(dff_q_5)
);
MUX2 mux_inst_1744 (
  .O(mux_o_1744),
  .I0(mux_o_1709),
  .I1(mux_o_1710),
  .S0(dff_q_5)
);
MUX2 mux_inst_1745 (
  .O(mux_o_1745),
  .I0(mux_o_1711),
  .I1(mux_o_1712),
  .S0(dff_q_5)
);
MUX2 mux_inst_1746 (
  .O(mux_o_1746),
  .I0(mux_o_1713),
  .I1(mux_o_1714),
  .S0(dff_q_5)
);
MUX2 mux_inst_1747 (
  .O(mux_o_1747),
  .I0(mux_o_1715),
  .I1(mux_o_1716),
  .S0(dff_q_4)
);
MUX2 mux_inst_1748 (
  .O(mux_o_1748),
  .I0(mux_o_1717),
  .I1(mux_o_1718),
  .S0(dff_q_4)
);
MUX2 mux_inst_1749 (
  .O(mux_o_1749),
  .I0(mux_o_1719),
  .I1(mux_o_1720),
  .S0(dff_q_4)
);
MUX2 mux_inst_1750 (
  .O(mux_o_1750),
  .I0(mux_o_1721),
  .I1(mux_o_1722),
  .S0(dff_q_4)
);
MUX2 mux_inst_1751 (
  .O(mux_o_1751),
  .I0(mux_o_1723),
  .I1(mux_o_1724),
  .S0(dff_q_4)
);
MUX2 mux_inst_1752 (
  .O(mux_o_1752),
  .I0(mux_o_1725),
  .I1(mux_o_1726),
  .S0(dff_q_4)
);
MUX2 mux_inst_1753 (
  .O(mux_o_1753),
  .I0(mux_o_1727),
  .I1(mux_o_1728),
  .S0(dff_q_4)
);
MUX2 mux_inst_1754 (
  .O(mux_o_1754),
  .I0(mux_o_1729),
  .I1(mux_o_1730),
  .S0(dff_q_4)
);
MUX2 mux_inst_1755 (
  .O(mux_o_1755),
  .I0(mux_o_1731),
  .I1(mux_o_1732),
  .S0(dff_q_4)
);
MUX2 mux_inst_1756 (
  .O(mux_o_1756),
  .I0(mux_o_1733),
  .I1(mux_o_1734),
  .S0(dff_q_4)
);
MUX2 mux_inst_1757 (
  .O(mux_o_1757),
  .I0(mux_o_1735),
  .I1(mux_o_1736),
  .S0(dff_q_4)
);
MUX2 mux_inst_1758 (
  .O(mux_o_1758),
  .I0(mux_o_1737),
  .I1(mux_o_1738),
  .S0(dff_q_4)
);
MUX2 mux_inst_1759 (
  .O(mux_o_1759),
  .I0(mux_o_1739),
  .I1(mux_o_1740),
  .S0(dff_q_4)
);
MUX2 mux_inst_1760 (
  .O(mux_o_1760),
  .I0(mux_o_1741),
  .I1(mux_o_1742),
  .S0(dff_q_4)
);
MUX2 mux_inst_1761 (
  .O(mux_o_1761),
  .I0(mux_o_1743),
  .I1(mux_o_1744),
  .S0(dff_q_4)
);
MUX2 mux_inst_1762 (
  .O(mux_o_1762),
  .I0(mux_o_1745),
  .I1(mux_o_1746),
  .S0(dff_q_4)
);
MUX2 mux_inst_1763 (
  .O(mux_o_1763),
  .I0(mux_o_1747),
  .I1(mux_o_1748),
  .S0(dff_q_3)
);
MUX2 mux_inst_1764 (
  .O(mux_o_1764),
  .I0(mux_o_1749),
  .I1(mux_o_1750),
  .S0(dff_q_3)
);
MUX2 mux_inst_1765 (
  .O(mux_o_1765),
  .I0(mux_o_1751),
  .I1(mux_o_1752),
  .S0(dff_q_3)
);
MUX2 mux_inst_1766 (
  .O(mux_o_1766),
  .I0(mux_o_1753),
  .I1(mux_o_1754),
  .S0(dff_q_3)
);
MUX2 mux_inst_1767 (
  .O(mux_o_1767),
  .I0(mux_o_1755),
  .I1(mux_o_1756),
  .S0(dff_q_3)
);
MUX2 mux_inst_1768 (
  .O(mux_o_1768),
  .I0(mux_o_1757),
  .I1(mux_o_1758),
  .S0(dff_q_3)
);
MUX2 mux_inst_1769 (
  .O(mux_o_1769),
  .I0(mux_o_1759),
  .I1(mux_o_1760),
  .S0(dff_q_3)
);
MUX2 mux_inst_1770 (
  .O(mux_o_1770),
  .I0(mux_o_1761),
  .I1(mux_o_1762),
  .S0(dff_q_3)
);
MUX2 mux_inst_1771 (
  .O(mux_o_1771),
  .I0(mux_o_1763),
  .I1(mux_o_1764),
  .S0(dff_q_2)
);
MUX2 mux_inst_1772 (
  .O(mux_o_1772),
  .I0(mux_o_1765),
  .I1(mux_o_1766),
  .S0(dff_q_2)
);
MUX2 mux_inst_1773 (
  .O(mux_o_1773),
  .I0(mux_o_1767),
  .I1(mux_o_1768),
  .S0(dff_q_2)
);
MUX2 mux_inst_1774 (
  .O(mux_o_1774),
  .I0(mux_o_1769),
  .I1(mux_o_1770),
  .S0(dff_q_2)
);
MUX2 mux_inst_1775 (
  .O(mux_o_1775),
  .I0(mux_o_1771),
  .I1(mux_o_1772),
  .S0(dff_q_1)
);
MUX2 mux_inst_1776 (
  .O(mux_o_1776),
  .I0(mux_o_1773),
  .I1(mux_o_1774),
  .S0(dff_q_1)
);
MUX2 mux_inst_1777 (
  .O(dout[13]),
  .I0(mux_o_1775),
  .I1(mux_o_1776),
  .S0(dff_q_0)
);
MUX2 mux_inst_1778 (
  .O(mux_o_1778),
  .I0(sdpb_inst_0_dout[14]),
  .I1(sdpb_inst_1_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1779 (
  .O(mux_o_1779),
  .I0(sdpb_inst_2_dout[14]),
  .I1(sdpb_inst_3_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1780 (
  .O(mux_o_1780),
  .I0(sdpb_inst_4_dout[14]),
  .I1(sdpb_inst_5_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1781 (
  .O(mux_o_1781),
  .I0(sdpb_inst_6_dout[14]),
  .I1(sdpb_inst_7_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1782 (
  .O(mux_o_1782),
  .I0(sdpb_inst_8_dout[14]),
  .I1(sdpb_inst_9_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1783 (
  .O(mux_o_1783),
  .I0(sdpb_inst_10_dout[14]),
  .I1(sdpb_inst_11_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1784 (
  .O(mux_o_1784),
  .I0(sdpb_inst_12_dout[14]),
  .I1(sdpb_inst_13_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1785 (
  .O(mux_o_1785),
  .I0(sdpb_inst_14_dout[14]),
  .I1(sdpb_inst_15_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1786 (
  .O(mux_o_1786),
  .I0(sdpb_inst_16_dout[14]),
  .I1(sdpb_inst_17_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1787 (
  .O(mux_o_1787),
  .I0(sdpb_inst_18_dout[14]),
  .I1(sdpb_inst_19_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1788 (
  .O(mux_o_1788),
  .I0(sdpb_inst_20_dout[14]),
  .I1(sdpb_inst_21_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1789 (
  .O(mux_o_1789),
  .I0(sdpb_inst_22_dout[14]),
  .I1(sdpb_inst_23_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1790 (
  .O(mux_o_1790),
  .I0(sdpb_inst_24_dout[14]),
  .I1(sdpb_inst_25_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1791 (
  .O(mux_o_1791),
  .I0(sdpb_inst_26_dout[14]),
  .I1(sdpb_inst_27_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1792 (
  .O(mux_o_1792),
  .I0(sdpb_inst_28_dout[14]),
  .I1(sdpb_inst_29_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1793 (
  .O(mux_o_1793),
  .I0(sdpb_inst_30_dout[14]),
  .I1(sdpb_inst_31_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1794 (
  .O(mux_o_1794),
  .I0(sdpb_inst_32_dout[14]),
  .I1(sdpb_inst_33_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1795 (
  .O(mux_o_1795),
  .I0(sdpb_inst_34_dout[14]),
  .I1(sdpb_inst_35_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1796 (
  .O(mux_o_1796),
  .I0(sdpb_inst_36_dout[14]),
  .I1(sdpb_inst_37_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1797 (
  .O(mux_o_1797),
  .I0(sdpb_inst_38_dout[14]),
  .I1(sdpb_inst_39_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1798 (
  .O(mux_o_1798),
  .I0(sdpb_inst_40_dout[14]),
  .I1(sdpb_inst_41_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1799 (
  .O(mux_o_1799),
  .I0(sdpb_inst_42_dout[14]),
  .I1(sdpb_inst_43_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1800 (
  .O(mux_o_1800),
  .I0(sdpb_inst_44_dout[14]),
  .I1(sdpb_inst_45_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1801 (
  .O(mux_o_1801),
  .I0(sdpb_inst_46_dout[14]),
  .I1(sdpb_inst_47_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1802 (
  .O(mux_o_1802),
  .I0(sdpb_inst_48_dout[14]),
  .I1(sdpb_inst_49_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1803 (
  .O(mux_o_1803),
  .I0(sdpb_inst_50_dout[14]),
  .I1(sdpb_inst_51_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1804 (
  .O(mux_o_1804),
  .I0(sdpb_inst_52_dout[14]),
  .I1(sdpb_inst_53_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1805 (
  .O(mux_o_1805),
  .I0(sdpb_inst_54_dout[14]),
  .I1(sdpb_inst_55_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1806 (
  .O(mux_o_1806),
  .I0(sdpb_inst_56_dout[14]),
  .I1(sdpb_inst_57_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1807 (
  .O(mux_o_1807),
  .I0(sdpb_inst_58_dout[14]),
  .I1(sdpb_inst_59_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1808 (
  .O(mux_o_1808),
  .I0(sdpb_inst_60_dout[14]),
  .I1(sdpb_inst_61_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1809 (
  .O(mux_o_1809),
  .I0(sdpb_inst_62_dout[14]),
  .I1(sdpb_inst_63_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1810 (
  .O(mux_o_1810),
  .I0(sdpb_inst_64_dout[14]),
  .I1(sdpb_inst_65_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1811 (
  .O(mux_o_1811),
  .I0(sdpb_inst_66_dout[14]),
  .I1(sdpb_inst_67_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1812 (
  .O(mux_o_1812),
  .I0(sdpb_inst_68_dout[14]),
  .I1(sdpb_inst_69_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1813 (
  .O(mux_o_1813),
  .I0(sdpb_inst_70_dout[14]),
  .I1(sdpb_inst_71_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1814 (
  .O(mux_o_1814),
  .I0(sdpb_inst_72_dout[14]),
  .I1(sdpb_inst_73_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1815 (
  .O(mux_o_1815),
  .I0(sdpb_inst_74_dout[14]),
  .I1(sdpb_inst_75_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1816 (
  .O(mux_o_1816),
  .I0(sdpb_inst_76_dout[14]),
  .I1(sdpb_inst_77_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1817 (
  .O(mux_o_1817),
  .I0(sdpb_inst_78_dout[14]),
  .I1(sdpb_inst_79_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1818 (
  .O(mux_o_1818),
  .I0(sdpb_inst_80_dout[14]),
  .I1(sdpb_inst_81_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1819 (
  .O(mux_o_1819),
  .I0(sdpb_inst_82_dout[14]),
  .I1(sdpb_inst_83_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1820 (
  .O(mux_o_1820),
  .I0(sdpb_inst_84_dout[14]),
  .I1(sdpb_inst_85_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1821 (
  .O(mux_o_1821),
  .I0(sdpb_inst_86_dout[14]),
  .I1(sdpb_inst_87_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1822 (
  .O(mux_o_1822),
  .I0(sdpb_inst_88_dout[14]),
  .I1(sdpb_inst_89_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1823 (
  .O(mux_o_1823),
  .I0(sdpb_inst_90_dout[14]),
  .I1(sdpb_inst_91_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1824 (
  .O(mux_o_1824),
  .I0(sdpb_inst_92_dout[14]),
  .I1(sdpb_inst_93_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1825 (
  .O(mux_o_1825),
  .I0(sdpb_inst_94_dout[14]),
  .I1(sdpb_inst_95_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1826 (
  .O(mux_o_1826),
  .I0(sdpb_inst_96_dout[14]),
  .I1(sdpb_inst_97_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1827 (
  .O(mux_o_1827),
  .I0(sdpb_inst_98_dout[14]),
  .I1(sdpb_inst_99_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1828 (
  .O(mux_o_1828),
  .I0(sdpb_inst_100_dout[14]),
  .I1(sdpb_inst_101_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1829 (
  .O(mux_o_1829),
  .I0(sdpb_inst_102_dout[14]),
  .I1(sdpb_inst_103_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1830 (
  .O(mux_o_1830),
  .I0(sdpb_inst_104_dout[14]),
  .I1(sdpb_inst_105_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1831 (
  .O(mux_o_1831),
  .I0(sdpb_inst_106_dout[14]),
  .I1(sdpb_inst_107_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1832 (
  .O(mux_o_1832),
  .I0(sdpb_inst_108_dout[14]),
  .I1(sdpb_inst_109_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1833 (
  .O(mux_o_1833),
  .I0(sdpb_inst_110_dout[14]),
  .I1(sdpb_inst_111_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1834 (
  .O(mux_o_1834),
  .I0(sdpb_inst_112_dout[14]),
  .I1(sdpb_inst_113_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1835 (
  .O(mux_o_1835),
  .I0(sdpb_inst_114_dout[14]),
  .I1(sdpb_inst_115_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1836 (
  .O(mux_o_1836),
  .I0(sdpb_inst_116_dout[14]),
  .I1(sdpb_inst_117_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1837 (
  .O(mux_o_1837),
  .I0(sdpb_inst_118_dout[14]),
  .I1(sdpb_inst_119_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1838 (
  .O(mux_o_1838),
  .I0(sdpb_inst_120_dout[14]),
  .I1(sdpb_inst_121_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1839 (
  .O(mux_o_1839),
  .I0(sdpb_inst_122_dout[14]),
  .I1(sdpb_inst_123_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1840 (
  .O(mux_o_1840),
  .I0(sdpb_inst_124_dout[14]),
  .I1(sdpb_inst_125_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1841 (
  .O(mux_o_1841),
  .I0(sdpb_inst_126_dout[14]),
  .I1(sdpb_inst_127_dout[14]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1842 (
  .O(mux_o_1842),
  .I0(mux_o_1778),
  .I1(mux_o_1779),
  .S0(dff_q_5)
);
MUX2 mux_inst_1843 (
  .O(mux_o_1843),
  .I0(mux_o_1780),
  .I1(mux_o_1781),
  .S0(dff_q_5)
);
MUX2 mux_inst_1844 (
  .O(mux_o_1844),
  .I0(mux_o_1782),
  .I1(mux_o_1783),
  .S0(dff_q_5)
);
MUX2 mux_inst_1845 (
  .O(mux_o_1845),
  .I0(mux_o_1784),
  .I1(mux_o_1785),
  .S0(dff_q_5)
);
MUX2 mux_inst_1846 (
  .O(mux_o_1846),
  .I0(mux_o_1786),
  .I1(mux_o_1787),
  .S0(dff_q_5)
);
MUX2 mux_inst_1847 (
  .O(mux_o_1847),
  .I0(mux_o_1788),
  .I1(mux_o_1789),
  .S0(dff_q_5)
);
MUX2 mux_inst_1848 (
  .O(mux_o_1848),
  .I0(mux_o_1790),
  .I1(mux_o_1791),
  .S0(dff_q_5)
);
MUX2 mux_inst_1849 (
  .O(mux_o_1849),
  .I0(mux_o_1792),
  .I1(mux_o_1793),
  .S0(dff_q_5)
);
MUX2 mux_inst_1850 (
  .O(mux_o_1850),
  .I0(mux_o_1794),
  .I1(mux_o_1795),
  .S0(dff_q_5)
);
MUX2 mux_inst_1851 (
  .O(mux_o_1851),
  .I0(mux_o_1796),
  .I1(mux_o_1797),
  .S0(dff_q_5)
);
MUX2 mux_inst_1852 (
  .O(mux_o_1852),
  .I0(mux_o_1798),
  .I1(mux_o_1799),
  .S0(dff_q_5)
);
MUX2 mux_inst_1853 (
  .O(mux_o_1853),
  .I0(mux_o_1800),
  .I1(mux_o_1801),
  .S0(dff_q_5)
);
MUX2 mux_inst_1854 (
  .O(mux_o_1854),
  .I0(mux_o_1802),
  .I1(mux_o_1803),
  .S0(dff_q_5)
);
MUX2 mux_inst_1855 (
  .O(mux_o_1855),
  .I0(mux_o_1804),
  .I1(mux_o_1805),
  .S0(dff_q_5)
);
MUX2 mux_inst_1856 (
  .O(mux_o_1856),
  .I0(mux_o_1806),
  .I1(mux_o_1807),
  .S0(dff_q_5)
);
MUX2 mux_inst_1857 (
  .O(mux_o_1857),
  .I0(mux_o_1808),
  .I1(mux_o_1809),
  .S0(dff_q_5)
);
MUX2 mux_inst_1858 (
  .O(mux_o_1858),
  .I0(mux_o_1810),
  .I1(mux_o_1811),
  .S0(dff_q_5)
);
MUX2 mux_inst_1859 (
  .O(mux_o_1859),
  .I0(mux_o_1812),
  .I1(mux_o_1813),
  .S0(dff_q_5)
);
MUX2 mux_inst_1860 (
  .O(mux_o_1860),
  .I0(mux_o_1814),
  .I1(mux_o_1815),
  .S0(dff_q_5)
);
MUX2 mux_inst_1861 (
  .O(mux_o_1861),
  .I0(mux_o_1816),
  .I1(mux_o_1817),
  .S0(dff_q_5)
);
MUX2 mux_inst_1862 (
  .O(mux_o_1862),
  .I0(mux_o_1818),
  .I1(mux_o_1819),
  .S0(dff_q_5)
);
MUX2 mux_inst_1863 (
  .O(mux_o_1863),
  .I0(mux_o_1820),
  .I1(mux_o_1821),
  .S0(dff_q_5)
);
MUX2 mux_inst_1864 (
  .O(mux_o_1864),
  .I0(mux_o_1822),
  .I1(mux_o_1823),
  .S0(dff_q_5)
);
MUX2 mux_inst_1865 (
  .O(mux_o_1865),
  .I0(mux_o_1824),
  .I1(mux_o_1825),
  .S0(dff_q_5)
);
MUX2 mux_inst_1866 (
  .O(mux_o_1866),
  .I0(mux_o_1826),
  .I1(mux_o_1827),
  .S0(dff_q_5)
);
MUX2 mux_inst_1867 (
  .O(mux_o_1867),
  .I0(mux_o_1828),
  .I1(mux_o_1829),
  .S0(dff_q_5)
);
MUX2 mux_inst_1868 (
  .O(mux_o_1868),
  .I0(mux_o_1830),
  .I1(mux_o_1831),
  .S0(dff_q_5)
);
MUX2 mux_inst_1869 (
  .O(mux_o_1869),
  .I0(mux_o_1832),
  .I1(mux_o_1833),
  .S0(dff_q_5)
);
MUX2 mux_inst_1870 (
  .O(mux_o_1870),
  .I0(mux_o_1834),
  .I1(mux_o_1835),
  .S0(dff_q_5)
);
MUX2 mux_inst_1871 (
  .O(mux_o_1871),
  .I0(mux_o_1836),
  .I1(mux_o_1837),
  .S0(dff_q_5)
);
MUX2 mux_inst_1872 (
  .O(mux_o_1872),
  .I0(mux_o_1838),
  .I1(mux_o_1839),
  .S0(dff_q_5)
);
MUX2 mux_inst_1873 (
  .O(mux_o_1873),
  .I0(mux_o_1840),
  .I1(mux_o_1841),
  .S0(dff_q_5)
);
MUX2 mux_inst_1874 (
  .O(mux_o_1874),
  .I0(mux_o_1842),
  .I1(mux_o_1843),
  .S0(dff_q_4)
);
MUX2 mux_inst_1875 (
  .O(mux_o_1875),
  .I0(mux_o_1844),
  .I1(mux_o_1845),
  .S0(dff_q_4)
);
MUX2 mux_inst_1876 (
  .O(mux_o_1876),
  .I0(mux_o_1846),
  .I1(mux_o_1847),
  .S0(dff_q_4)
);
MUX2 mux_inst_1877 (
  .O(mux_o_1877),
  .I0(mux_o_1848),
  .I1(mux_o_1849),
  .S0(dff_q_4)
);
MUX2 mux_inst_1878 (
  .O(mux_o_1878),
  .I0(mux_o_1850),
  .I1(mux_o_1851),
  .S0(dff_q_4)
);
MUX2 mux_inst_1879 (
  .O(mux_o_1879),
  .I0(mux_o_1852),
  .I1(mux_o_1853),
  .S0(dff_q_4)
);
MUX2 mux_inst_1880 (
  .O(mux_o_1880),
  .I0(mux_o_1854),
  .I1(mux_o_1855),
  .S0(dff_q_4)
);
MUX2 mux_inst_1881 (
  .O(mux_o_1881),
  .I0(mux_o_1856),
  .I1(mux_o_1857),
  .S0(dff_q_4)
);
MUX2 mux_inst_1882 (
  .O(mux_o_1882),
  .I0(mux_o_1858),
  .I1(mux_o_1859),
  .S0(dff_q_4)
);
MUX2 mux_inst_1883 (
  .O(mux_o_1883),
  .I0(mux_o_1860),
  .I1(mux_o_1861),
  .S0(dff_q_4)
);
MUX2 mux_inst_1884 (
  .O(mux_o_1884),
  .I0(mux_o_1862),
  .I1(mux_o_1863),
  .S0(dff_q_4)
);
MUX2 mux_inst_1885 (
  .O(mux_o_1885),
  .I0(mux_o_1864),
  .I1(mux_o_1865),
  .S0(dff_q_4)
);
MUX2 mux_inst_1886 (
  .O(mux_o_1886),
  .I0(mux_o_1866),
  .I1(mux_o_1867),
  .S0(dff_q_4)
);
MUX2 mux_inst_1887 (
  .O(mux_o_1887),
  .I0(mux_o_1868),
  .I1(mux_o_1869),
  .S0(dff_q_4)
);
MUX2 mux_inst_1888 (
  .O(mux_o_1888),
  .I0(mux_o_1870),
  .I1(mux_o_1871),
  .S0(dff_q_4)
);
MUX2 mux_inst_1889 (
  .O(mux_o_1889),
  .I0(mux_o_1872),
  .I1(mux_o_1873),
  .S0(dff_q_4)
);
MUX2 mux_inst_1890 (
  .O(mux_o_1890),
  .I0(mux_o_1874),
  .I1(mux_o_1875),
  .S0(dff_q_3)
);
MUX2 mux_inst_1891 (
  .O(mux_o_1891),
  .I0(mux_o_1876),
  .I1(mux_o_1877),
  .S0(dff_q_3)
);
MUX2 mux_inst_1892 (
  .O(mux_o_1892),
  .I0(mux_o_1878),
  .I1(mux_o_1879),
  .S0(dff_q_3)
);
MUX2 mux_inst_1893 (
  .O(mux_o_1893),
  .I0(mux_o_1880),
  .I1(mux_o_1881),
  .S0(dff_q_3)
);
MUX2 mux_inst_1894 (
  .O(mux_o_1894),
  .I0(mux_o_1882),
  .I1(mux_o_1883),
  .S0(dff_q_3)
);
MUX2 mux_inst_1895 (
  .O(mux_o_1895),
  .I0(mux_o_1884),
  .I1(mux_o_1885),
  .S0(dff_q_3)
);
MUX2 mux_inst_1896 (
  .O(mux_o_1896),
  .I0(mux_o_1886),
  .I1(mux_o_1887),
  .S0(dff_q_3)
);
MUX2 mux_inst_1897 (
  .O(mux_o_1897),
  .I0(mux_o_1888),
  .I1(mux_o_1889),
  .S0(dff_q_3)
);
MUX2 mux_inst_1898 (
  .O(mux_o_1898),
  .I0(mux_o_1890),
  .I1(mux_o_1891),
  .S0(dff_q_2)
);
MUX2 mux_inst_1899 (
  .O(mux_o_1899),
  .I0(mux_o_1892),
  .I1(mux_o_1893),
  .S0(dff_q_2)
);
MUX2 mux_inst_1900 (
  .O(mux_o_1900),
  .I0(mux_o_1894),
  .I1(mux_o_1895),
  .S0(dff_q_2)
);
MUX2 mux_inst_1901 (
  .O(mux_o_1901),
  .I0(mux_o_1896),
  .I1(mux_o_1897),
  .S0(dff_q_2)
);
MUX2 mux_inst_1902 (
  .O(mux_o_1902),
  .I0(mux_o_1898),
  .I1(mux_o_1899),
  .S0(dff_q_1)
);
MUX2 mux_inst_1903 (
  .O(mux_o_1903),
  .I0(mux_o_1900),
  .I1(mux_o_1901),
  .S0(dff_q_1)
);
MUX2 mux_inst_1904 (
  .O(dout[14]),
  .I0(mux_o_1902),
  .I1(mux_o_1903),
  .S0(dff_q_0)
);
MUX2 mux_inst_1905 (
  .O(mux_o_1905),
  .I0(sdpb_inst_0_dout[15]),
  .I1(sdpb_inst_1_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1906 (
  .O(mux_o_1906),
  .I0(sdpb_inst_2_dout[15]),
  .I1(sdpb_inst_3_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1907 (
  .O(mux_o_1907),
  .I0(sdpb_inst_4_dout[15]),
  .I1(sdpb_inst_5_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1908 (
  .O(mux_o_1908),
  .I0(sdpb_inst_6_dout[15]),
  .I1(sdpb_inst_7_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1909 (
  .O(mux_o_1909),
  .I0(sdpb_inst_8_dout[15]),
  .I1(sdpb_inst_9_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1910 (
  .O(mux_o_1910),
  .I0(sdpb_inst_10_dout[15]),
  .I1(sdpb_inst_11_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1911 (
  .O(mux_o_1911),
  .I0(sdpb_inst_12_dout[15]),
  .I1(sdpb_inst_13_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1912 (
  .O(mux_o_1912),
  .I0(sdpb_inst_14_dout[15]),
  .I1(sdpb_inst_15_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1913 (
  .O(mux_o_1913),
  .I0(sdpb_inst_16_dout[15]),
  .I1(sdpb_inst_17_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1914 (
  .O(mux_o_1914),
  .I0(sdpb_inst_18_dout[15]),
  .I1(sdpb_inst_19_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1915 (
  .O(mux_o_1915),
  .I0(sdpb_inst_20_dout[15]),
  .I1(sdpb_inst_21_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1916 (
  .O(mux_o_1916),
  .I0(sdpb_inst_22_dout[15]),
  .I1(sdpb_inst_23_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1917 (
  .O(mux_o_1917),
  .I0(sdpb_inst_24_dout[15]),
  .I1(sdpb_inst_25_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1918 (
  .O(mux_o_1918),
  .I0(sdpb_inst_26_dout[15]),
  .I1(sdpb_inst_27_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1919 (
  .O(mux_o_1919),
  .I0(sdpb_inst_28_dout[15]),
  .I1(sdpb_inst_29_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1920 (
  .O(mux_o_1920),
  .I0(sdpb_inst_30_dout[15]),
  .I1(sdpb_inst_31_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1921 (
  .O(mux_o_1921),
  .I0(sdpb_inst_32_dout[15]),
  .I1(sdpb_inst_33_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1922 (
  .O(mux_o_1922),
  .I0(sdpb_inst_34_dout[15]),
  .I1(sdpb_inst_35_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1923 (
  .O(mux_o_1923),
  .I0(sdpb_inst_36_dout[15]),
  .I1(sdpb_inst_37_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1924 (
  .O(mux_o_1924),
  .I0(sdpb_inst_38_dout[15]),
  .I1(sdpb_inst_39_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1925 (
  .O(mux_o_1925),
  .I0(sdpb_inst_40_dout[15]),
  .I1(sdpb_inst_41_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1926 (
  .O(mux_o_1926),
  .I0(sdpb_inst_42_dout[15]),
  .I1(sdpb_inst_43_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1927 (
  .O(mux_o_1927),
  .I0(sdpb_inst_44_dout[15]),
  .I1(sdpb_inst_45_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1928 (
  .O(mux_o_1928),
  .I0(sdpb_inst_46_dout[15]),
  .I1(sdpb_inst_47_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1929 (
  .O(mux_o_1929),
  .I0(sdpb_inst_48_dout[15]),
  .I1(sdpb_inst_49_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1930 (
  .O(mux_o_1930),
  .I0(sdpb_inst_50_dout[15]),
  .I1(sdpb_inst_51_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1931 (
  .O(mux_o_1931),
  .I0(sdpb_inst_52_dout[15]),
  .I1(sdpb_inst_53_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1932 (
  .O(mux_o_1932),
  .I0(sdpb_inst_54_dout[15]),
  .I1(sdpb_inst_55_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1933 (
  .O(mux_o_1933),
  .I0(sdpb_inst_56_dout[15]),
  .I1(sdpb_inst_57_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1934 (
  .O(mux_o_1934),
  .I0(sdpb_inst_58_dout[15]),
  .I1(sdpb_inst_59_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1935 (
  .O(mux_o_1935),
  .I0(sdpb_inst_60_dout[15]),
  .I1(sdpb_inst_61_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1936 (
  .O(mux_o_1936),
  .I0(sdpb_inst_62_dout[15]),
  .I1(sdpb_inst_63_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1937 (
  .O(mux_o_1937),
  .I0(sdpb_inst_64_dout[15]),
  .I1(sdpb_inst_65_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1938 (
  .O(mux_o_1938),
  .I0(sdpb_inst_66_dout[15]),
  .I1(sdpb_inst_67_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1939 (
  .O(mux_o_1939),
  .I0(sdpb_inst_68_dout[15]),
  .I1(sdpb_inst_69_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1940 (
  .O(mux_o_1940),
  .I0(sdpb_inst_70_dout[15]),
  .I1(sdpb_inst_71_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1941 (
  .O(mux_o_1941),
  .I0(sdpb_inst_72_dout[15]),
  .I1(sdpb_inst_73_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1942 (
  .O(mux_o_1942),
  .I0(sdpb_inst_74_dout[15]),
  .I1(sdpb_inst_75_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1943 (
  .O(mux_o_1943),
  .I0(sdpb_inst_76_dout[15]),
  .I1(sdpb_inst_77_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1944 (
  .O(mux_o_1944),
  .I0(sdpb_inst_78_dout[15]),
  .I1(sdpb_inst_79_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1945 (
  .O(mux_o_1945),
  .I0(sdpb_inst_80_dout[15]),
  .I1(sdpb_inst_81_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1946 (
  .O(mux_o_1946),
  .I0(sdpb_inst_82_dout[15]),
  .I1(sdpb_inst_83_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1947 (
  .O(mux_o_1947),
  .I0(sdpb_inst_84_dout[15]),
  .I1(sdpb_inst_85_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1948 (
  .O(mux_o_1948),
  .I0(sdpb_inst_86_dout[15]),
  .I1(sdpb_inst_87_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1949 (
  .O(mux_o_1949),
  .I0(sdpb_inst_88_dout[15]),
  .I1(sdpb_inst_89_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1950 (
  .O(mux_o_1950),
  .I0(sdpb_inst_90_dout[15]),
  .I1(sdpb_inst_91_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1951 (
  .O(mux_o_1951),
  .I0(sdpb_inst_92_dout[15]),
  .I1(sdpb_inst_93_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1952 (
  .O(mux_o_1952),
  .I0(sdpb_inst_94_dout[15]),
  .I1(sdpb_inst_95_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1953 (
  .O(mux_o_1953),
  .I0(sdpb_inst_96_dout[15]),
  .I1(sdpb_inst_97_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1954 (
  .O(mux_o_1954),
  .I0(sdpb_inst_98_dout[15]),
  .I1(sdpb_inst_99_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1955 (
  .O(mux_o_1955),
  .I0(sdpb_inst_100_dout[15]),
  .I1(sdpb_inst_101_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1956 (
  .O(mux_o_1956),
  .I0(sdpb_inst_102_dout[15]),
  .I1(sdpb_inst_103_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1957 (
  .O(mux_o_1957),
  .I0(sdpb_inst_104_dout[15]),
  .I1(sdpb_inst_105_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1958 (
  .O(mux_o_1958),
  .I0(sdpb_inst_106_dout[15]),
  .I1(sdpb_inst_107_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1959 (
  .O(mux_o_1959),
  .I0(sdpb_inst_108_dout[15]),
  .I1(sdpb_inst_109_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1960 (
  .O(mux_o_1960),
  .I0(sdpb_inst_110_dout[15]),
  .I1(sdpb_inst_111_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1961 (
  .O(mux_o_1961),
  .I0(sdpb_inst_112_dout[15]),
  .I1(sdpb_inst_113_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1962 (
  .O(mux_o_1962),
  .I0(sdpb_inst_114_dout[15]),
  .I1(sdpb_inst_115_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1963 (
  .O(mux_o_1963),
  .I0(sdpb_inst_116_dout[15]),
  .I1(sdpb_inst_117_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1964 (
  .O(mux_o_1964),
  .I0(sdpb_inst_118_dout[15]),
  .I1(sdpb_inst_119_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1965 (
  .O(mux_o_1965),
  .I0(sdpb_inst_120_dout[15]),
  .I1(sdpb_inst_121_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1966 (
  .O(mux_o_1966),
  .I0(sdpb_inst_122_dout[15]),
  .I1(sdpb_inst_123_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1967 (
  .O(mux_o_1967),
  .I0(sdpb_inst_124_dout[15]),
  .I1(sdpb_inst_125_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1968 (
  .O(mux_o_1968),
  .I0(sdpb_inst_126_dout[15]),
  .I1(sdpb_inst_127_dout[15]),
  .S0(dff_q_6)
);
MUX2 mux_inst_1969 (
  .O(mux_o_1969),
  .I0(mux_o_1905),
  .I1(mux_o_1906),
  .S0(dff_q_5)
);
MUX2 mux_inst_1970 (
  .O(mux_o_1970),
  .I0(mux_o_1907),
  .I1(mux_o_1908),
  .S0(dff_q_5)
);
MUX2 mux_inst_1971 (
  .O(mux_o_1971),
  .I0(mux_o_1909),
  .I1(mux_o_1910),
  .S0(dff_q_5)
);
MUX2 mux_inst_1972 (
  .O(mux_o_1972),
  .I0(mux_o_1911),
  .I1(mux_o_1912),
  .S0(dff_q_5)
);
MUX2 mux_inst_1973 (
  .O(mux_o_1973),
  .I0(mux_o_1913),
  .I1(mux_o_1914),
  .S0(dff_q_5)
);
MUX2 mux_inst_1974 (
  .O(mux_o_1974),
  .I0(mux_o_1915),
  .I1(mux_o_1916),
  .S0(dff_q_5)
);
MUX2 mux_inst_1975 (
  .O(mux_o_1975),
  .I0(mux_o_1917),
  .I1(mux_o_1918),
  .S0(dff_q_5)
);
MUX2 mux_inst_1976 (
  .O(mux_o_1976),
  .I0(mux_o_1919),
  .I1(mux_o_1920),
  .S0(dff_q_5)
);
MUX2 mux_inst_1977 (
  .O(mux_o_1977),
  .I0(mux_o_1921),
  .I1(mux_o_1922),
  .S0(dff_q_5)
);
MUX2 mux_inst_1978 (
  .O(mux_o_1978),
  .I0(mux_o_1923),
  .I1(mux_o_1924),
  .S0(dff_q_5)
);
MUX2 mux_inst_1979 (
  .O(mux_o_1979),
  .I0(mux_o_1925),
  .I1(mux_o_1926),
  .S0(dff_q_5)
);
MUX2 mux_inst_1980 (
  .O(mux_o_1980),
  .I0(mux_o_1927),
  .I1(mux_o_1928),
  .S0(dff_q_5)
);
MUX2 mux_inst_1981 (
  .O(mux_o_1981),
  .I0(mux_o_1929),
  .I1(mux_o_1930),
  .S0(dff_q_5)
);
MUX2 mux_inst_1982 (
  .O(mux_o_1982),
  .I0(mux_o_1931),
  .I1(mux_o_1932),
  .S0(dff_q_5)
);
MUX2 mux_inst_1983 (
  .O(mux_o_1983),
  .I0(mux_o_1933),
  .I1(mux_o_1934),
  .S0(dff_q_5)
);
MUX2 mux_inst_1984 (
  .O(mux_o_1984),
  .I0(mux_o_1935),
  .I1(mux_o_1936),
  .S0(dff_q_5)
);
MUX2 mux_inst_1985 (
  .O(mux_o_1985),
  .I0(mux_o_1937),
  .I1(mux_o_1938),
  .S0(dff_q_5)
);
MUX2 mux_inst_1986 (
  .O(mux_o_1986),
  .I0(mux_o_1939),
  .I1(mux_o_1940),
  .S0(dff_q_5)
);
MUX2 mux_inst_1987 (
  .O(mux_o_1987),
  .I0(mux_o_1941),
  .I1(mux_o_1942),
  .S0(dff_q_5)
);
MUX2 mux_inst_1988 (
  .O(mux_o_1988),
  .I0(mux_o_1943),
  .I1(mux_o_1944),
  .S0(dff_q_5)
);
MUX2 mux_inst_1989 (
  .O(mux_o_1989),
  .I0(mux_o_1945),
  .I1(mux_o_1946),
  .S0(dff_q_5)
);
MUX2 mux_inst_1990 (
  .O(mux_o_1990),
  .I0(mux_o_1947),
  .I1(mux_o_1948),
  .S0(dff_q_5)
);
MUX2 mux_inst_1991 (
  .O(mux_o_1991),
  .I0(mux_o_1949),
  .I1(mux_o_1950),
  .S0(dff_q_5)
);
MUX2 mux_inst_1992 (
  .O(mux_o_1992),
  .I0(mux_o_1951),
  .I1(mux_o_1952),
  .S0(dff_q_5)
);
MUX2 mux_inst_1993 (
  .O(mux_o_1993),
  .I0(mux_o_1953),
  .I1(mux_o_1954),
  .S0(dff_q_5)
);
MUX2 mux_inst_1994 (
  .O(mux_o_1994),
  .I0(mux_o_1955),
  .I1(mux_o_1956),
  .S0(dff_q_5)
);
MUX2 mux_inst_1995 (
  .O(mux_o_1995),
  .I0(mux_o_1957),
  .I1(mux_o_1958),
  .S0(dff_q_5)
);
MUX2 mux_inst_1996 (
  .O(mux_o_1996),
  .I0(mux_o_1959),
  .I1(mux_o_1960),
  .S0(dff_q_5)
);
MUX2 mux_inst_1997 (
  .O(mux_o_1997),
  .I0(mux_o_1961),
  .I1(mux_o_1962),
  .S0(dff_q_5)
);
MUX2 mux_inst_1998 (
  .O(mux_o_1998),
  .I0(mux_o_1963),
  .I1(mux_o_1964),
  .S0(dff_q_5)
);
MUX2 mux_inst_1999 (
  .O(mux_o_1999),
  .I0(mux_o_1965),
  .I1(mux_o_1966),
  .S0(dff_q_5)
);
MUX2 mux_inst_2000 (
  .O(mux_o_2000),
  .I0(mux_o_1967),
  .I1(mux_o_1968),
  .S0(dff_q_5)
);
MUX2 mux_inst_2001 (
  .O(mux_o_2001),
  .I0(mux_o_1969),
  .I1(mux_o_1970),
  .S0(dff_q_4)
);
MUX2 mux_inst_2002 (
  .O(mux_o_2002),
  .I0(mux_o_1971),
  .I1(mux_o_1972),
  .S0(dff_q_4)
);
MUX2 mux_inst_2003 (
  .O(mux_o_2003),
  .I0(mux_o_1973),
  .I1(mux_o_1974),
  .S0(dff_q_4)
);
MUX2 mux_inst_2004 (
  .O(mux_o_2004),
  .I0(mux_o_1975),
  .I1(mux_o_1976),
  .S0(dff_q_4)
);
MUX2 mux_inst_2005 (
  .O(mux_o_2005),
  .I0(mux_o_1977),
  .I1(mux_o_1978),
  .S0(dff_q_4)
);
MUX2 mux_inst_2006 (
  .O(mux_o_2006),
  .I0(mux_o_1979),
  .I1(mux_o_1980),
  .S0(dff_q_4)
);
MUX2 mux_inst_2007 (
  .O(mux_o_2007),
  .I0(mux_o_1981),
  .I1(mux_o_1982),
  .S0(dff_q_4)
);
MUX2 mux_inst_2008 (
  .O(mux_o_2008),
  .I0(mux_o_1983),
  .I1(mux_o_1984),
  .S0(dff_q_4)
);
MUX2 mux_inst_2009 (
  .O(mux_o_2009),
  .I0(mux_o_1985),
  .I1(mux_o_1986),
  .S0(dff_q_4)
);
MUX2 mux_inst_2010 (
  .O(mux_o_2010),
  .I0(mux_o_1987),
  .I1(mux_o_1988),
  .S0(dff_q_4)
);
MUX2 mux_inst_2011 (
  .O(mux_o_2011),
  .I0(mux_o_1989),
  .I1(mux_o_1990),
  .S0(dff_q_4)
);
MUX2 mux_inst_2012 (
  .O(mux_o_2012),
  .I0(mux_o_1991),
  .I1(mux_o_1992),
  .S0(dff_q_4)
);
MUX2 mux_inst_2013 (
  .O(mux_o_2013),
  .I0(mux_o_1993),
  .I1(mux_o_1994),
  .S0(dff_q_4)
);
MUX2 mux_inst_2014 (
  .O(mux_o_2014),
  .I0(mux_o_1995),
  .I1(mux_o_1996),
  .S0(dff_q_4)
);
MUX2 mux_inst_2015 (
  .O(mux_o_2015),
  .I0(mux_o_1997),
  .I1(mux_o_1998),
  .S0(dff_q_4)
);
MUX2 mux_inst_2016 (
  .O(mux_o_2016),
  .I0(mux_o_1999),
  .I1(mux_o_2000),
  .S0(dff_q_4)
);
MUX2 mux_inst_2017 (
  .O(mux_o_2017),
  .I0(mux_o_2001),
  .I1(mux_o_2002),
  .S0(dff_q_3)
);
MUX2 mux_inst_2018 (
  .O(mux_o_2018),
  .I0(mux_o_2003),
  .I1(mux_o_2004),
  .S0(dff_q_3)
);
MUX2 mux_inst_2019 (
  .O(mux_o_2019),
  .I0(mux_o_2005),
  .I1(mux_o_2006),
  .S0(dff_q_3)
);
MUX2 mux_inst_2020 (
  .O(mux_o_2020),
  .I0(mux_o_2007),
  .I1(mux_o_2008),
  .S0(dff_q_3)
);
MUX2 mux_inst_2021 (
  .O(mux_o_2021),
  .I0(mux_o_2009),
  .I1(mux_o_2010),
  .S0(dff_q_3)
);
MUX2 mux_inst_2022 (
  .O(mux_o_2022),
  .I0(mux_o_2011),
  .I1(mux_o_2012),
  .S0(dff_q_3)
);
MUX2 mux_inst_2023 (
  .O(mux_o_2023),
  .I0(mux_o_2013),
  .I1(mux_o_2014),
  .S0(dff_q_3)
);
MUX2 mux_inst_2024 (
  .O(mux_o_2024),
  .I0(mux_o_2015),
  .I1(mux_o_2016),
  .S0(dff_q_3)
);
MUX2 mux_inst_2025 (
  .O(mux_o_2025),
  .I0(mux_o_2017),
  .I1(mux_o_2018),
  .S0(dff_q_2)
);
MUX2 mux_inst_2026 (
  .O(mux_o_2026),
  .I0(mux_o_2019),
  .I1(mux_o_2020),
  .S0(dff_q_2)
);
MUX2 mux_inst_2027 (
  .O(mux_o_2027),
  .I0(mux_o_2021),
  .I1(mux_o_2022),
  .S0(dff_q_2)
);
MUX2 mux_inst_2028 (
  .O(mux_o_2028),
  .I0(mux_o_2023),
  .I1(mux_o_2024),
  .S0(dff_q_2)
);
MUX2 mux_inst_2029 (
  .O(mux_o_2029),
  .I0(mux_o_2025),
  .I1(mux_o_2026),
  .S0(dff_q_1)
);
MUX2 mux_inst_2030 (
  .O(mux_o_2030),
  .I0(mux_o_2027),
  .I1(mux_o_2028),
  .S0(dff_q_1)
);
MUX2 mux_inst_2031 (
  .O(dout[15]),
  .I0(mux_o_2029),
  .I1(mux_o_2030),
  .S0(dff_q_0)
);
MUX2 mux_inst_2032 (
  .O(mux_o_2032),
  .I0(sdpb_inst_128_dout[16]),
  .I1(sdpb_inst_129_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2033 (
  .O(mux_o_2033),
  .I0(sdpb_inst_130_dout[16]),
  .I1(sdpb_inst_131_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2034 (
  .O(mux_o_2034),
  .I0(sdpb_inst_132_dout[16]),
  .I1(sdpb_inst_133_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2035 (
  .O(mux_o_2035),
  .I0(sdpb_inst_134_dout[16]),
  .I1(sdpb_inst_135_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2036 (
  .O(mux_o_2036),
  .I0(sdpb_inst_136_dout[16]),
  .I1(sdpb_inst_137_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2037 (
  .O(mux_o_2037),
  .I0(sdpb_inst_138_dout[16]),
  .I1(sdpb_inst_139_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2038 (
  .O(mux_o_2038),
  .I0(sdpb_inst_140_dout[16]),
  .I1(sdpb_inst_141_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2039 (
  .O(mux_o_2039),
  .I0(sdpb_inst_142_dout[16]),
  .I1(sdpb_inst_143_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2040 (
  .O(mux_o_2040),
  .I0(sdpb_inst_144_dout[16]),
  .I1(sdpb_inst_145_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2041 (
  .O(mux_o_2041),
  .I0(sdpb_inst_146_dout[16]),
  .I1(sdpb_inst_147_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2042 (
  .O(mux_o_2042),
  .I0(sdpb_inst_148_dout[16]),
  .I1(sdpb_inst_149_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2043 (
  .O(mux_o_2043),
  .I0(sdpb_inst_150_dout[16]),
  .I1(sdpb_inst_151_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2044 (
  .O(mux_o_2044),
  .I0(sdpb_inst_152_dout[16]),
  .I1(sdpb_inst_153_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2045 (
  .O(mux_o_2045),
  .I0(sdpb_inst_154_dout[16]),
  .I1(sdpb_inst_155_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2046 (
  .O(mux_o_2046),
  .I0(sdpb_inst_156_dout[16]),
  .I1(sdpb_inst_157_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2047 (
  .O(mux_o_2047),
  .I0(sdpb_inst_158_dout[16]),
  .I1(sdpb_inst_159_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2048 (
  .O(mux_o_2048),
  .I0(sdpb_inst_160_dout[16]),
  .I1(sdpb_inst_161_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2049 (
  .O(mux_o_2049),
  .I0(sdpb_inst_162_dout[16]),
  .I1(sdpb_inst_163_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2050 (
  .O(mux_o_2050),
  .I0(sdpb_inst_164_dout[16]),
  .I1(sdpb_inst_165_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2051 (
  .O(mux_o_2051),
  .I0(sdpb_inst_166_dout[16]),
  .I1(sdpb_inst_167_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2052 (
  .O(mux_o_2052),
  .I0(sdpb_inst_168_dout[16]),
  .I1(sdpb_inst_169_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2053 (
  .O(mux_o_2053),
  .I0(sdpb_inst_170_dout[16]),
  .I1(sdpb_inst_171_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2054 (
  .O(mux_o_2054),
  .I0(sdpb_inst_172_dout[16]),
  .I1(sdpb_inst_173_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2055 (
  .O(mux_o_2055),
  .I0(sdpb_inst_174_dout[16]),
  .I1(sdpb_inst_175_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2056 (
  .O(mux_o_2056),
  .I0(sdpb_inst_176_dout[16]),
  .I1(sdpb_inst_177_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2057 (
  .O(mux_o_2057),
  .I0(sdpb_inst_178_dout[16]),
  .I1(sdpb_inst_179_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2058 (
  .O(mux_o_2058),
  .I0(sdpb_inst_180_dout[16]),
  .I1(sdpb_inst_181_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2059 (
  .O(mux_o_2059),
  .I0(sdpb_inst_182_dout[16]),
  .I1(sdpb_inst_183_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2060 (
  .O(mux_o_2060),
  .I0(sdpb_inst_184_dout[16]),
  .I1(sdpb_inst_185_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2061 (
  .O(mux_o_2061),
  .I0(sdpb_inst_186_dout[16]),
  .I1(sdpb_inst_187_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2062 (
  .O(mux_o_2062),
  .I0(sdpb_inst_188_dout[16]),
  .I1(sdpb_inst_189_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2063 (
  .O(mux_o_2063),
  .I0(sdpb_inst_190_dout[16]),
  .I1(sdpb_inst_191_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2064 (
  .O(mux_o_2064),
  .I0(sdpb_inst_192_dout[16]),
  .I1(sdpb_inst_193_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2065 (
  .O(mux_o_2065),
  .I0(sdpb_inst_194_dout[16]),
  .I1(sdpb_inst_195_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2066 (
  .O(mux_o_2066),
  .I0(sdpb_inst_196_dout[16]),
  .I1(sdpb_inst_197_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2067 (
  .O(mux_o_2067),
  .I0(sdpb_inst_198_dout[16]),
  .I1(sdpb_inst_199_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2068 (
  .O(mux_o_2068),
  .I0(sdpb_inst_200_dout[16]),
  .I1(sdpb_inst_201_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2069 (
  .O(mux_o_2069),
  .I0(sdpb_inst_202_dout[16]),
  .I1(sdpb_inst_203_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2070 (
  .O(mux_o_2070),
  .I0(sdpb_inst_204_dout[16]),
  .I1(sdpb_inst_205_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2071 (
  .O(mux_o_2071),
  .I0(sdpb_inst_206_dout[16]),
  .I1(sdpb_inst_207_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2072 (
  .O(mux_o_2072),
  .I0(sdpb_inst_208_dout[16]),
  .I1(sdpb_inst_209_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2073 (
  .O(mux_o_2073),
  .I0(sdpb_inst_210_dout[16]),
  .I1(sdpb_inst_211_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2074 (
  .O(mux_o_2074),
  .I0(sdpb_inst_212_dout[16]),
  .I1(sdpb_inst_213_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2075 (
  .O(mux_o_2075),
  .I0(sdpb_inst_214_dout[16]),
  .I1(sdpb_inst_215_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2076 (
  .O(mux_o_2076),
  .I0(sdpb_inst_216_dout[16]),
  .I1(sdpb_inst_217_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2077 (
  .O(mux_o_2077),
  .I0(sdpb_inst_218_dout[16]),
  .I1(sdpb_inst_219_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2078 (
  .O(mux_o_2078),
  .I0(sdpb_inst_220_dout[16]),
  .I1(sdpb_inst_221_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2079 (
  .O(mux_o_2079),
  .I0(sdpb_inst_222_dout[16]),
  .I1(sdpb_inst_223_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2080 (
  .O(mux_o_2080),
  .I0(sdpb_inst_224_dout[16]),
  .I1(sdpb_inst_225_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2081 (
  .O(mux_o_2081),
  .I0(sdpb_inst_226_dout[16]),
  .I1(sdpb_inst_227_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2082 (
  .O(mux_o_2082),
  .I0(sdpb_inst_228_dout[16]),
  .I1(sdpb_inst_229_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2083 (
  .O(mux_o_2083),
  .I0(sdpb_inst_230_dout[16]),
  .I1(sdpb_inst_231_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2084 (
  .O(mux_o_2084),
  .I0(sdpb_inst_232_dout[16]),
  .I1(sdpb_inst_233_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2085 (
  .O(mux_o_2085),
  .I0(sdpb_inst_234_dout[16]),
  .I1(sdpb_inst_235_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2086 (
  .O(mux_o_2086),
  .I0(sdpb_inst_236_dout[16]),
  .I1(sdpb_inst_237_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2087 (
  .O(mux_o_2087),
  .I0(sdpb_inst_238_dout[16]),
  .I1(sdpb_inst_239_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2088 (
  .O(mux_o_2088),
  .I0(sdpb_inst_240_dout[16]),
  .I1(sdpb_inst_241_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2089 (
  .O(mux_o_2089),
  .I0(sdpb_inst_242_dout[16]),
  .I1(sdpb_inst_243_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2090 (
  .O(mux_o_2090),
  .I0(sdpb_inst_244_dout[16]),
  .I1(sdpb_inst_245_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2091 (
  .O(mux_o_2091),
  .I0(sdpb_inst_246_dout[16]),
  .I1(sdpb_inst_247_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2092 (
  .O(mux_o_2092),
  .I0(sdpb_inst_248_dout[16]),
  .I1(sdpb_inst_249_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2093 (
  .O(mux_o_2093),
  .I0(sdpb_inst_250_dout[16]),
  .I1(sdpb_inst_251_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2094 (
  .O(mux_o_2094),
  .I0(sdpb_inst_252_dout[16]),
  .I1(sdpb_inst_253_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2095 (
  .O(mux_o_2095),
  .I0(sdpb_inst_254_dout[16]),
  .I1(sdpb_inst_255_dout[16]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2096 (
  .O(mux_o_2096),
  .I0(mux_o_2032),
  .I1(mux_o_2033),
  .S0(dff_q_5)
);
MUX2 mux_inst_2097 (
  .O(mux_o_2097),
  .I0(mux_o_2034),
  .I1(mux_o_2035),
  .S0(dff_q_5)
);
MUX2 mux_inst_2098 (
  .O(mux_o_2098),
  .I0(mux_o_2036),
  .I1(mux_o_2037),
  .S0(dff_q_5)
);
MUX2 mux_inst_2099 (
  .O(mux_o_2099),
  .I0(mux_o_2038),
  .I1(mux_o_2039),
  .S0(dff_q_5)
);
MUX2 mux_inst_2100 (
  .O(mux_o_2100),
  .I0(mux_o_2040),
  .I1(mux_o_2041),
  .S0(dff_q_5)
);
MUX2 mux_inst_2101 (
  .O(mux_o_2101),
  .I0(mux_o_2042),
  .I1(mux_o_2043),
  .S0(dff_q_5)
);
MUX2 mux_inst_2102 (
  .O(mux_o_2102),
  .I0(mux_o_2044),
  .I1(mux_o_2045),
  .S0(dff_q_5)
);
MUX2 mux_inst_2103 (
  .O(mux_o_2103),
  .I0(mux_o_2046),
  .I1(mux_o_2047),
  .S0(dff_q_5)
);
MUX2 mux_inst_2104 (
  .O(mux_o_2104),
  .I0(mux_o_2048),
  .I1(mux_o_2049),
  .S0(dff_q_5)
);
MUX2 mux_inst_2105 (
  .O(mux_o_2105),
  .I0(mux_o_2050),
  .I1(mux_o_2051),
  .S0(dff_q_5)
);
MUX2 mux_inst_2106 (
  .O(mux_o_2106),
  .I0(mux_o_2052),
  .I1(mux_o_2053),
  .S0(dff_q_5)
);
MUX2 mux_inst_2107 (
  .O(mux_o_2107),
  .I0(mux_o_2054),
  .I1(mux_o_2055),
  .S0(dff_q_5)
);
MUX2 mux_inst_2108 (
  .O(mux_o_2108),
  .I0(mux_o_2056),
  .I1(mux_o_2057),
  .S0(dff_q_5)
);
MUX2 mux_inst_2109 (
  .O(mux_o_2109),
  .I0(mux_o_2058),
  .I1(mux_o_2059),
  .S0(dff_q_5)
);
MUX2 mux_inst_2110 (
  .O(mux_o_2110),
  .I0(mux_o_2060),
  .I1(mux_o_2061),
  .S0(dff_q_5)
);
MUX2 mux_inst_2111 (
  .O(mux_o_2111),
  .I0(mux_o_2062),
  .I1(mux_o_2063),
  .S0(dff_q_5)
);
MUX2 mux_inst_2112 (
  .O(mux_o_2112),
  .I0(mux_o_2064),
  .I1(mux_o_2065),
  .S0(dff_q_5)
);
MUX2 mux_inst_2113 (
  .O(mux_o_2113),
  .I0(mux_o_2066),
  .I1(mux_o_2067),
  .S0(dff_q_5)
);
MUX2 mux_inst_2114 (
  .O(mux_o_2114),
  .I0(mux_o_2068),
  .I1(mux_o_2069),
  .S0(dff_q_5)
);
MUX2 mux_inst_2115 (
  .O(mux_o_2115),
  .I0(mux_o_2070),
  .I1(mux_o_2071),
  .S0(dff_q_5)
);
MUX2 mux_inst_2116 (
  .O(mux_o_2116),
  .I0(mux_o_2072),
  .I1(mux_o_2073),
  .S0(dff_q_5)
);
MUX2 mux_inst_2117 (
  .O(mux_o_2117),
  .I0(mux_o_2074),
  .I1(mux_o_2075),
  .S0(dff_q_5)
);
MUX2 mux_inst_2118 (
  .O(mux_o_2118),
  .I0(mux_o_2076),
  .I1(mux_o_2077),
  .S0(dff_q_5)
);
MUX2 mux_inst_2119 (
  .O(mux_o_2119),
  .I0(mux_o_2078),
  .I1(mux_o_2079),
  .S0(dff_q_5)
);
MUX2 mux_inst_2120 (
  .O(mux_o_2120),
  .I0(mux_o_2080),
  .I1(mux_o_2081),
  .S0(dff_q_5)
);
MUX2 mux_inst_2121 (
  .O(mux_o_2121),
  .I0(mux_o_2082),
  .I1(mux_o_2083),
  .S0(dff_q_5)
);
MUX2 mux_inst_2122 (
  .O(mux_o_2122),
  .I0(mux_o_2084),
  .I1(mux_o_2085),
  .S0(dff_q_5)
);
MUX2 mux_inst_2123 (
  .O(mux_o_2123),
  .I0(mux_o_2086),
  .I1(mux_o_2087),
  .S0(dff_q_5)
);
MUX2 mux_inst_2124 (
  .O(mux_o_2124),
  .I0(mux_o_2088),
  .I1(mux_o_2089),
  .S0(dff_q_5)
);
MUX2 mux_inst_2125 (
  .O(mux_o_2125),
  .I0(mux_o_2090),
  .I1(mux_o_2091),
  .S0(dff_q_5)
);
MUX2 mux_inst_2126 (
  .O(mux_o_2126),
  .I0(mux_o_2092),
  .I1(mux_o_2093),
  .S0(dff_q_5)
);
MUX2 mux_inst_2127 (
  .O(mux_o_2127),
  .I0(mux_o_2094),
  .I1(mux_o_2095),
  .S0(dff_q_5)
);
MUX2 mux_inst_2128 (
  .O(mux_o_2128),
  .I0(mux_o_2096),
  .I1(mux_o_2097),
  .S0(dff_q_4)
);
MUX2 mux_inst_2129 (
  .O(mux_o_2129),
  .I0(mux_o_2098),
  .I1(mux_o_2099),
  .S0(dff_q_4)
);
MUX2 mux_inst_2130 (
  .O(mux_o_2130),
  .I0(mux_o_2100),
  .I1(mux_o_2101),
  .S0(dff_q_4)
);
MUX2 mux_inst_2131 (
  .O(mux_o_2131),
  .I0(mux_o_2102),
  .I1(mux_o_2103),
  .S0(dff_q_4)
);
MUX2 mux_inst_2132 (
  .O(mux_o_2132),
  .I0(mux_o_2104),
  .I1(mux_o_2105),
  .S0(dff_q_4)
);
MUX2 mux_inst_2133 (
  .O(mux_o_2133),
  .I0(mux_o_2106),
  .I1(mux_o_2107),
  .S0(dff_q_4)
);
MUX2 mux_inst_2134 (
  .O(mux_o_2134),
  .I0(mux_o_2108),
  .I1(mux_o_2109),
  .S0(dff_q_4)
);
MUX2 mux_inst_2135 (
  .O(mux_o_2135),
  .I0(mux_o_2110),
  .I1(mux_o_2111),
  .S0(dff_q_4)
);
MUX2 mux_inst_2136 (
  .O(mux_o_2136),
  .I0(mux_o_2112),
  .I1(mux_o_2113),
  .S0(dff_q_4)
);
MUX2 mux_inst_2137 (
  .O(mux_o_2137),
  .I0(mux_o_2114),
  .I1(mux_o_2115),
  .S0(dff_q_4)
);
MUX2 mux_inst_2138 (
  .O(mux_o_2138),
  .I0(mux_o_2116),
  .I1(mux_o_2117),
  .S0(dff_q_4)
);
MUX2 mux_inst_2139 (
  .O(mux_o_2139),
  .I0(mux_o_2118),
  .I1(mux_o_2119),
  .S0(dff_q_4)
);
MUX2 mux_inst_2140 (
  .O(mux_o_2140),
  .I0(mux_o_2120),
  .I1(mux_o_2121),
  .S0(dff_q_4)
);
MUX2 mux_inst_2141 (
  .O(mux_o_2141),
  .I0(mux_o_2122),
  .I1(mux_o_2123),
  .S0(dff_q_4)
);
MUX2 mux_inst_2142 (
  .O(mux_o_2142),
  .I0(mux_o_2124),
  .I1(mux_o_2125),
  .S0(dff_q_4)
);
MUX2 mux_inst_2143 (
  .O(mux_o_2143),
  .I0(mux_o_2126),
  .I1(mux_o_2127),
  .S0(dff_q_4)
);
MUX2 mux_inst_2144 (
  .O(mux_o_2144),
  .I0(mux_o_2128),
  .I1(mux_o_2129),
  .S0(dff_q_3)
);
MUX2 mux_inst_2145 (
  .O(mux_o_2145),
  .I0(mux_o_2130),
  .I1(mux_o_2131),
  .S0(dff_q_3)
);
MUX2 mux_inst_2146 (
  .O(mux_o_2146),
  .I0(mux_o_2132),
  .I1(mux_o_2133),
  .S0(dff_q_3)
);
MUX2 mux_inst_2147 (
  .O(mux_o_2147),
  .I0(mux_o_2134),
  .I1(mux_o_2135),
  .S0(dff_q_3)
);
MUX2 mux_inst_2148 (
  .O(mux_o_2148),
  .I0(mux_o_2136),
  .I1(mux_o_2137),
  .S0(dff_q_3)
);
MUX2 mux_inst_2149 (
  .O(mux_o_2149),
  .I0(mux_o_2138),
  .I1(mux_o_2139),
  .S0(dff_q_3)
);
MUX2 mux_inst_2150 (
  .O(mux_o_2150),
  .I0(mux_o_2140),
  .I1(mux_o_2141),
  .S0(dff_q_3)
);
MUX2 mux_inst_2151 (
  .O(mux_o_2151),
  .I0(mux_o_2142),
  .I1(mux_o_2143),
  .S0(dff_q_3)
);
MUX2 mux_inst_2152 (
  .O(mux_o_2152),
  .I0(mux_o_2144),
  .I1(mux_o_2145),
  .S0(dff_q_2)
);
MUX2 mux_inst_2153 (
  .O(mux_o_2153),
  .I0(mux_o_2146),
  .I1(mux_o_2147),
  .S0(dff_q_2)
);
MUX2 mux_inst_2154 (
  .O(mux_o_2154),
  .I0(mux_o_2148),
  .I1(mux_o_2149),
  .S0(dff_q_2)
);
MUX2 mux_inst_2155 (
  .O(mux_o_2155),
  .I0(mux_o_2150),
  .I1(mux_o_2151),
  .S0(dff_q_2)
);
MUX2 mux_inst_2156 (
  .O(mux_o_2156),
  .I0(mux_o_2152),
  .I1(mux_o_2153),
  .S0(dff_q_1)
);
MUX2 mux_inst_2157 (
  .O(mux_o_2157),
  .I0(mux_o_2154),
  .I1(mux_o_2155),
  .S0(dff_q_1)
);
MUX2 mux_inst_2158 (
  .O(dout[16]),
  .I0(mux_o_2156),
  .I1(mux_o_2157),
  .S0(dff_q_0)
);
MUX2 mux_inst_2159 (
  .O(mux_o_2159),
  .I0(sdpb_inst_128_dout[17]),
  .I1(sdpb_inst_129_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2160 (
  .O(mux_o_2160),
  .I0(sdpb_inst_130_dout[17]),
  .I1(sdpb_inst_131_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2161 (
  .O(mux_o_2161),
  .I0(sdpb_inst_132_dout[17]),
  .I1(sdpb_inst_133_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2162 (
  .O(mux_o_2162),
  .I0(sdpb_inst_134_dout[17]),
  .I1(sdpb_inst_135_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2163 (
  .O(mux_o_2163),
  .I0(sdpb_inst_136_dout[17]),
  .I1(sdpb_inst_137_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2164 (
  .O(mux_o_2164),
  .I0(sdpb_inst_138_dout[17]),
  .I1(sdpb_inst_139_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2165 (
  .O(mux_o_2165),
  .I0(sdpb_inst_140_dout[17]),
  .I1(sdpb_inst_141_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2166 (
  .O(mux_o_2166),
  .I0(sdpb_inst_142_dout[17]),
  .I1(sdpb_inst_143_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2167 (
  .O(mux_o_2167),
  .I0(sdpb_inst_144_dout[17]),
  .I1(sdpb_inst_145_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2168 (
  .O(mux_o_2168),
  .I0(sdpb_inst_146_dout[17]),
  .I1(sdpb_inst_147_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2169 (
  .O(mux_o_2169),
  .I0(sdpb_inst_148_dout[17]),
  .I1(sdpb_inst_149_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2170 (
  .O(mux_o_2170),
  .I0(sdpb_inst_150_dout[17]),
  .I1(sdpb_inst_151_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2171 (
  .O(mux_o_2171),
  .I0(sdpb_inst_152_dout[17]),
  .I1(sdpb_inst_153_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2172 (
  .O(mux_o_2172),
  .I0(sdpb_inst_154_dout[17]),
  .I1(sdpb_inst_155_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2173 (
  .O(mux_o_2173),
  .I0(sdpb_inst_156_dout[17]),
  .I1(sdpb_inst_157_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2174 (
  .O(mux_o_2174),
  .I0(sdpb_inst_158_dout[17]),
  .I1(sdpb_inst_159_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2175 (
  .O(mux_o_2175),
  .I0(sdpb_inst_160_dout[17]),
  .I1(sdpb_inst_161_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2176 (
  .O(mux_o_2176),
  .I0(sdpb_inst_162_dout[17]),
  .I1(sdpb_inst_163_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2177 (
  .O(mux_o_2177),
  .I0(sdpb_inst_164_dout[17]),
  .I1(sdpb_inst_165_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2178 (
  .O(mux_o_2178),
  .I0(sdpb_inst_166_dout[17]),
  .I1(sdpb_inst_167_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2179 (
  .O(mux_o_2179),
  .I0(sdpb_inst_168_dout[17]),
  .I1(sdpb_inst_169_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2180 (
  .O(mux_o_2180),
  .I0(sdpb_inst_170_dout[17]),
  .I1(sdpb_inst_171_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2181 (
  .O(mux_o_2181),
  .I0(sdpb_inst_172_dout[17]),
  .I1(sdpb_inst_173_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2182 (
  .O(mux_o_2182),
  .I0(sdpb_inst_174_dout[17]),
  .I1(sdpb_inst_175_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2183 (
  .O(mux_o_2183),
  .I0(sdpb_inst_176_dout[17]),
  .I1(sdpb_inst_177_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2184 (
  .O(mux_o_2184),
  .I0(sdpb_inst_178_dout[17]),
  .I1(sdpb_inst_179_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2185 (
  .O(mux_o_2185),
  .I0(sdpb_inst_180_dout[17]),
  .I1(sdpb_inst_181_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2186 (
  .O(mux_o_2186),
  .I0(sdpb_inst_182_dout[17]),
  .I1(sdpb_inst_183_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2187 (
  .O(mux_o_2187),
  .I0(sdpb_inst_184_dout[17]),
  .I1(sdpb_inst_185_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2188 (
  .O(mux_o_2188),
  .I0(sdpb_inst_186_dout[17]),
  .I1(sdpb_inst_187_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2189 (
  .O(mux_o_2189),
  .I0(sdpb_inst_188_dout[17]),
  .I1(sdpb_inst_189_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2190 (
  .O(mux_o_2190),
  .I0(sdpb_inst_190_dout[17]),
  .I1(sdpb_inst_191_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2191 (
  .O(mux_o_2191),
  .I0(sdpb_inst_192_dout[17]),
  .I1(sdpb_inst_193_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2192 (
  .O(mux_o_2192),
  .I0(sdpb_inst_194_dout[17]),
  .I1(sdpb_inst_195_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2193 (
  .O(mux_o_2193),
  .I0(sdpb_inst_196_dout[17]),
  .I1(sdpb_inst_197_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2194 (
  .O(mux_o_2194),
  .I0(sdpb_inst_198_dout[17]),
  .I1(sdpb_inst_199_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2195 (
  .O(mux_o_2195),
  .I0(sdpb_inst_200_dout[17]),
  .I1(sdpb_inst_201_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2196 (
  .O(mux_o_2196),
  .I0(sdpb_inst_202_dout[17]),
  .I1(sdpb_inst_203_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2197 (
  .O(mux_o_2197),
  .I0(sdpb_inst_204_dout[17]),
  .I1(sdpb_inst_205_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2198 (
  .O(mux_o_2198),
  .I0(sdpb_inst_206_dout[17]),
  .I1(sdpb_inst_207_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2199 (
  .O(mux_o_2199),
  .I0(sdpb_inst_208_dout[17]),
  .I1(sdpb_inst_209_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2200 (
  .O(mux_o_2200),
  .I0(sdpb_inst_210_dout[17]),
  .I1(sdpb_inst_211_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2201 (
  .O(mux_o_2201),
  .I0(sdpb_inst_212_dout[17]),
  .I1(sdpb_inst_213_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2202 (
  .O(mux_o_2202),
  .I0(sdpb_inst_214_dout[17]),
  .I1(sdpb_inst_215_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2203 (
  .O(mux_o_2203),
  .I0(sdpb_inst_216_dout[17]),
  .I1(sdpb_inst_217_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2204 (
  .O(mux_o_2204),
  .I0(sdpb_inst_218_dout[17]),
  .I1(sdpb_inst_219_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2205 (
  .O(mux_o_2205),
  .I0(sdpb_inst_220_dout[17]),
  .I1(sdpb_inst_221_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2206 (
  .O(mux_o_2206),
  .I0(sdpb_inst_222_dout[17]),
  .I1(sdpb_inst_223_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2207 (
  .O(mux_o_2207),
  .I0(sdpb_inst_224_dout[17]),
  .I1(sdpb_inst_225_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2208 (
  .O(mux_o_2208),
  .I0(sdpb_inst_226_dout[17]),
  .I1(sdpb_inst_227_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2209 (
  .O(mux_o_2209),
  .I0(sdpb_inst_228_dout[17]),
  .I1(sdpb_inst_229_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2210 (
  .O(mux_o_2210),
  .I0(sdpb_inst_230_dout[17]),
  .I1(sdpb_inst_231_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2211 (
  .O(mux_o_2211),
  .I0(sdpb_inst_232_dout[17]),
  .I1(sdpb_inst_233_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2212 (
  .O(mux_o_2212),
  .I0(sdpb_inst_234_dout[17]),
  .I1(sdpb_inst_235_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2213 (
  .O(mux_o_2213),
  .I0(sdpb_inst_236_dout[17]),
  .I1(sdpb_inst_237_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2214 (
  .O(mux_o_2214),
  .I0(sdpb_inst_238_dout[17]),
  .I1(sdpb_inst_239_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2215 (
  .O(mux_o_2215),
  .I0(sdpb_inst_240_dout[17]),
  .I1(sdpb_inst_241_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2216 (
  .O(mux_o_2216),
  .I0(sdpb_inst_242_dout[17]),
  .I1(sdpb_inst_243_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2217 (
  .O(mux_o_2217),
  .I0(sdpb_inst_244_dout[17]),
  .I1(sdpb_inst_245_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2218 (
  .O(mux_o_2218),
  .I0(sdpb_inst_246_dout[17]),
  .I1(sdpb_inst_247_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2219 (
  .O(mux_o_2219),
  .I0(sdpb_inst_248_dout[17]),
  .I1(sdpb_inst_249_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2220 (
  .O(mux_o_2220),
  .I0(sdpb_inst_250_dout[17]),
  .I1(sdpb_inst_251_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2221 (
  .O(mux_o_2221),
  .I0(sdpb_inst_252_dout[17]),
  .I1(sdpb_inst_253_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2222 (
  .O(mux_o_2222),
  .I0(sdpb_inst_254_dout[17]),
  .I1(sdpb_inst_255_dout[17]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2223 (
  .O(mux_o_2223),
  .I0(mux_o_2159),
  .I1(mux_o_2160),
  .S0(dff_q_5)
);
MUX2 mux_inst_2224 (
  .O(mux_o_2224),
  .I0(mux_o_2161),
  .I1(mux_o_2162),
  .S0(dff_q_5)
);
MUX2 mux_inst_2225 (
  .O(mux_o_2225),
  .I0(mux_o_2163),
  .I1(mux_o_2164),
  .S0(dff_q_5)
);
MUX2 mux_inst_2226 (
  .O(mux_o_2226),
  .I0(mux_o_2165),
  .I1(mux_o_2166),
  .S0(dff_q_5)
);
MUX2 mux_inst_2227 (
  .O(mux_o_2227),
  .I0(mux_o_2167),
  .I1(mux_o_2168),
  .S0(dff_q_5)
);
MUX2 mux_inst_2228 (
  .O(mux_o_2228),
  .I0(mux_o_2169),
  .I1(mux_o_2170),
  .S0(dff_q_5)
);
MUX2 mux_inst_2229 (
  .O(mux_o_2229),
  .I0(mux_o_2171),
  .I1(mux_o_2172),
  .S0(dff_q_5)
);
MUX2 mux_inst_2230 (
  .O(mux_o_2230),
  .I0(mux_o_2173),
  .I1(mux_o_2174),
  .S0(dff_q_5)
);
MUX2 mux_inst_2231 (
  .O(mux_o_2231),
  .I0(mux_o_2175),
  .I1(mux_o_2176),
  .S0(dff_q_5)
);
MUX2 mux_inst_2232 (
  .O(mux_o_2232),
  .I0(mux_o_2177),
  .I1(mux_o_2178),
  .S0(dff_q_5)
);
MUX2 mux_inst_2233 (
  .O(mux_o_2233),
  .I0(mux_o_2179),
  .I1(mux_o_2180),
  .S0(dff_q_5)
);
MUX2 mux_inst_2234 (
  .O(mux_o_2234),
  .I0(mux_o_2181),
  .I1(mux_o_2182),
  .S0(dff_q_5)
);
MUX2 mux_inst_2235 (
  .O(mux_o_2235),
  .I0(mux_o_2183),
  .I1(mux_o_2184),
  .S0(dff_q_5)
);
MUX2 mux_inst_2236 (
  .O(mux_o_2236),
  .I0(mux_o_2185),
  .I1(mux_o_2186),
  .S0(dff_q_5)
);
MUX2 mux_inst_2237 (
  .O(mux_o_2237),
  .I0(mux_o_2187),
  .I1(mux_o_2188),
  .S0(dff_q_5)
);
MUX2 mux_inst_2238 (
  .O(mux_o_2238),
  .I0(mux_o_2189),
  .I1(mux_o_2190),
  .S0(dff_q_5)
);
MUX2 mux_inst_2239 (
  .O(mux_o_2239),
  .I0(mux_o_2191),
  .I1(mux_o_2192),
  .S0(dff_q_5)
);
MUX2 mux_inst_2240 (
  .O(mux_o_2240),
  .I0(mux_o_2193),
  .I1(mux_o_2194),
  .S0(dff_q_5)
);
MUX2 mux_inst_2241 (
  .O(mux_o_2241),
  .I0(mux_o_2195),
  .I1(mux_o_2196),
  .S0(dff_q_5)
);
MUX2 mux_inst_2242 (
  .O(mux_o_2242),
  .I0(mux_o_2197),
  .I1(mux_o_2198),
  .S0(dff_q_5)
);
MUX2 mux_inst_2243 (
  .O(mux_o_2243),
  .I0(mux_o_2199),
  .I1(mux_o_2200),
  .S0(dff_q_5)
);
MUX2 mux_inst_2244 (
  .O(mux_o_2244),
  .I0(mux_o_2201),
  .I1(mux_o_2202),
  .S0(dff_q_5)
);
MUX2 mux_inst_2245 (
  .O(mux_o_2245),
  .I0(mux_o_2203),
  .I1(mux_o_2204),
  .S0(dff_q_5)
);
MUX2 mux_inst_2246 (
  .O(mux_o_2246),
  .I0(mux_o_2205),
  .I1(mux_o_2206),
  .S0(dff_q_5)
);
MUX2 mux_inst_2247 (
  .O(mux_o_2247),
  .I0(mux_o_2207),
  .I1(mux_o_2208),
  .S0(dff_q_5)
);
MUX2 mux_inst_2248 (
  .O(mux_o_2248),
  .I0(mux_o_2209),
  .I1(mux_o_2210),
  .S0(dff_q_5)
);
MUX2 mux_inst_2249 (
  .O(mux_o_2249),
  .I0(mux_o_2211),
  .I1(mux_o_2212),
  .S0(dff_q_5)
);
MUX2 mux_inst_2250 (
  .O(mux_o_2250),
  .I0(mux_o_2213),
  .I1(mux_o_2214),
  .S0(dff_q_5)
);
MUX2 mux_inst_2251 (
  .O(mux_o_2251),
  .I0(mux_o_2215),
  .I1(mux_o_2216),
  .S0(dff_q_5)
);
MUX2 mux_inst_2252 (
  .O(mux_o_2252),
  .I0(mux_o_2217),
  .I1(mux_o_2218),
  .S0(dff_q_5)
);
MUX2 mux_inst_2253 (
  .O(mux_o_2253),
  .I0(mux_o_2219),
  .I1(mux_o_2220),
  .S0(dff_q_5)
);
MUX2 mux_inst_2254 (
  .O(mux_o_2254),
  .I0(mux_o_2221),
  .I1(mux_o_2222),
  .S0(dff_q_5)
);
MUX2 mux_inst_2255 (
  .O(mux_o_2255),
  .I0(mux_o_2223),
  .I1(mux_o_2224),
  .S0(dff_q_4)
);
MUX2 mux_inst_2256 (
  .O(mux_o_2256),
  .I0(mux_o_2225),
  .I1(mux_o_2226),
  .S0(dff_q_4)
);
MUX2 mux_inst_2257 (
  .O(mux_o_2257),
  .I0(mux_o_2227),
  .I1(mux_o_2228),
  .S0(dff_q_4)
);
MUX2 mux_inst_2258 (
  .O(mux_o_2258),
  .I0(mux_o_2229),
  .I1(mux_o_2230),
  .S0(dff_q_4)
);
MUX2 mux_inst_2259 (
  .O(mux_o_2259),
  .I0(mux_o_2231),
  .I1(mux_o_2232),
  .S0(dff_q_4)
);
MUX2 mux_inst_2260 (
  .O(mux_o_2260),
  .I0(mux_o_2233),
  .I1(mux_o_2234),
  .S0(dff_q_4)
);
MUX2 mux_inst_2261 (
  .O(mux_o_2261),
  .I0(mux_o_2235),
  .I1(mux_o_2236),
  .S0(dff_q_4)
);
MUX2 mux_inst_2262 (
  .O(mux_o_2262),
  .I0(mux_o_2237),
  .I1(mux_o_2238),
  .S0(dff_q_4)
);
MUX2 mux_inst_2263 (
  .O(mux_o_2263),
  .I0(mux_o_2239),
  .I1(mux_o_2240),
  .S0(dff_q_4)
);
MUX2 mux_inst_2264 (
  .O(mux_o_2264),
  .I0(mux_o_2241),
  .I1(mux_o_2242),
  .S0(dff_q_4)
);
MUX2 mux_inst_2265 (
  .O(mux_o_2265),
  .I0(mux_o_2243),
  .I1(mux_o_2244),
  .S0(dff_q_4)
);
MUX2 mux_inst_2266 (
  .O(mux_o_2266),
  .I0(mux_o_2245),
  .I1(mux_o_2246),
  .S0(dff_q_4)
);
MUX2 mux_inst_2267 (
  .O(mux_o_2267),
  .I0(mux_o_2247),
  .I1(mux_o_2248),
  .S0(dff_q_4)
);
MUX2 mux_inst_2268 (
  .O(mux_o_2268),
  .I0(mux_o_2249),
  .I1(mux_o_2250),
  .S0(dff_q_4)
);
MUX2 mux_inst_2269 (
  .O(mux_o_2269),
  .I0(mux_o_2251),
  .I1(mux_o_2252),
  .S0(dff_q_4)
);
MUX2 mux_inst_2270 (
  .O(mux_o_2270),
  .I0(mux_o_2253),
  .I1(mux_o_2254),
  .S0(dff_q_4)
);
MUX2 mux_inst_2271 (
  .O(mux_o_2271),
  .I0(mux_o_2255),
  .I1(mux_o_2256),
  .S0(dff_q_3)
);
MUX2 mux_inst_2272 (
  .O(mux_o_2272),
  .I0(mux_o_2257),
  .I1(mux_o_2258),
  .S0(dff_q_3)
);
MUX2 mux_inst_2273 (
  .O(mux_o_2273),
  .I0(mux_o_2259),
  .I1(mux_o_2260),
  .S0(dff_q_3)
);
MUX2 mux_inst_2274 (
  .O(mux_o_2274),
  .I0(mux_o_2261),
  .I1(mux_o_2262),
  .S0(dff_q_3)
);
MUX2 mux_inst_2275 (
  .O(mux_o_2275),
  .I0(mux_o_2263),
  .I1(mux_o_2264),
  .S0(dff_q_3)
);
MUX2 mux_inst_2276 (
  .O(mux_o_2276),
  .I0(mux_o_2265),
  .I1(mux_o_2266),
  .S0(dff_q_3)
);
MUX2 mux_inst_2277 (
  .O(mux_o_2277),
  .I0(mux_o_2267),
  .I1(mux_o_2268),
  .S0(dff_q_3)
);
MUX2 mux_inst_2278 (
  .O(mux_o_2278),
  .I0(mux_o_2269),
  .I1(mux_o_2270),
  .S0(dff_q_3)
);
MUX2 mux_inst_2279 (
  .O(mux_o_2279),
  .I0(mux_o_2271),
  .I1(mux_o_2272),
  .S0(dff_q_2)
);
MUX2 mux_inst_2280 (
  .O(mux_o_2280),
  .I0(mux_o_2273),
  .I1(mux_o_2274),
  .S0(dff_q_2)
);
MUX2 mux_inst_2281 (
  .O(mux_o_2281),
  .I0(mux_o_2275),
  .I1(mux_o_2276),
  .S0(dff_q_2)
);
MUX2 mux_inst_2282 (
  .O(mux_o_2282),
  .I0(mux_o_2277),
  .I1(mux_o_2278),
  .S0(dff_q_2)
);
MUX2 mux_inst_2283 (
  .O(mux_o_2283),
  .I0(mux_o_2279),
  .I1(mux_o_2280),
  .S0(dff_q_1)
);
MUX2 mux_inst_2284 (
  .O(mux_o_2284),
  .I0(mux_o_2281),
  .I1(mux_o_2282),
  .S0(dff_q_1)
);
MUX2 mux_inst_2285 (
  .O(dout[17]),
  .I0(mux_o_2283),
  .I1(mux_o_2284),
  .S0(dff_q_0)
);
MUX2 mux_inst_2286 (
  .O(mux_o_2286),
  .I0(sdpb_inst_128_dout[18]),
  .I1(sdpb_inst_129_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2287 (
  .O(mux_o_2287),
  .I0(sdpb_inst_130_dout[18]),
  .I1(sdpb_inst_131_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2288 (
  .O(mux_o_2288),
  .I0(sdpb_inst_132_dout[18]),
  .I1(sdpb_inst_133_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2289 (
  .O(mux_o_2289),
  .I0(sdpb_inst_134_dout[18]),
  .I1(sdpb_inst_135_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2290 (
  .O(mux_o_2290),
  .I0(sdpb_inst_136_dout[18]),
  .I1(sdpb_inst_137_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2291 (
  .O(mux_o_2291),
  .I0(sdpb_inst_138_dout[18]),
  .I1(sdpb_inst_139_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2292 (
  .O(mux_o_2292),
  .I0(sdpb_inst_140_dout[18]),
  .I1(sdpb_inst_141_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2293 (
  .O(mux_o_2293),
  .I0(sdpb_inst_142_dout[18]),
  .I1(sdpb_inst_143_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2294 (
  .O(mux_o_2294),
  .I0(sdpb_inst_144_dout[18]),
  .I1(sdpb_inst_145_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2295 (
  .O(mux_o_2295),
  .I0(sdpb_inst_146_dout[18]),
  .I1(sdpb_inst_147_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2296 (
  .O(mux_o_2296),
  .I0(sdpb_inst_148_dout[18]),
  .I1(sdpb_inst_149_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2297 (
  .O(mux_o_2297),
  .I0(sdpb_inst_150_dout[18]),
  .I1(sdpb_inst_151_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2298 (
  .O(mux_o_2298),
  .I0(sdpb_inst_152_dout[18]),
  .I1(sdpb_inst_153_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2299 (
  .O(mux_o_2299),
  .I0(sdpb_inst_154_dout[18]),
  .I1(sdpb_inst_155_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2300 (
  .O(mux_o_2300),
  .I0(sdpb_inst_156_dout[18]),
  .I1(sdpb_inst_157_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2301 (
  .O(mux_o_2301),
  .I0(sdpb_inst_158_dout[18]),
  .I1(sdpb_inst_159_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2302 (
  .O(mux_o_2302),
  .I0(sdpb_inst_160_dout[18]),
  .I1(sdpb_inst_161_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2303 (
  .O(mux_o_2303),
  .I0(sdpb_inst_162_dout[18]),
  .I1(sdpb_inst_163_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2304 (
  .O(mux_o_2304),
  .I0(sdpb_inst_164_dout[18]),
  .I1(sdpb_inst_165_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2305 (
  .O(mux_o_2305),
  .I0(sdpb_inst_166_dout[18]),
  .I1(sdpb_inst_167_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2306 (
  .O(mux_o_2306),
  .I0(sdpb_inst_168_dout[18]),
  .I1(sdpb_inst_169_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2307 (
  .O(mux_o_2307),
  .I0(sdpb_inst_170_dout[18]),
  .I1(sdpb_inst_171_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2308 (
  .O(mux_o_2308),
  .I0(sdpb_inst_172_dout[18]),
  .I1(sdpb_inst_173_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2309 (
  .O(mux_o_2309),
  .I0(sdpb_inst_174_dout[18]),
  .I1(sdpb_inst_175_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2310 (
  .O(mux_o_2310),
  .I0(sdpb_inst_176_dout[18]),
  .I1(sdpb_inst_177_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2311 (
  .O(mux_o_2311),
  .I0(sdpb_inst_178_dout[18]),
  .I1(sdpb_inst_179_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2312 (
  .O(mux_o_2312),
  .I0(sdpb_inst_180_dout[18]),
  .I1(sdpb_inst_181_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2313 (
  .O(mux_o_2313),
  .I0(sdpb_inst_182_dout[18]),
  .I1(sdpb_inst_183_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2314 (
  .O(mux_o_2314),
  .I0(sdpb_inst_184_dout[18]),
  .I1(sdpb_inst_185_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2315 (
  .O(mux_o_2315),
  .I0(sdpb_inst_186_dout[18]),
  .I1(sdpb_inst_187_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2316 (
  .O(mux_o_2316),
  .I0(sdpb_inst_188_dout[18]),
  .I1(sdpb_inst_189_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2317 (
  .O(mux_o_2317),
  .I0(sdpb_inst_190_dout[18]),
  .I1(sdpb_inst_191_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2318 (
  .O(mux_o_2318),
  .I0(sdpb_inst_192_dout[18]),
  .I1(sdpb_inst_193_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2319 (
  .O(mux_o_2319),
  .I0(sdpb_inst_194_dout[18]),
  .I1(sdpb_inst_195_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2320 (
  .O(mux_o_2320),
  .I0(sdpb_inst_196_dout[18]),
  .I1(sdpb_inst_197_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2321 (
  .O(mux_o_2321),
  .I0(sdpb_inst_198_dout[18]),
  .I1(sdpb_inst_199_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2322 (
  .O(mux_o_2322),
  .I0(sdpb_inst_200_dout[18]),
  .I1(sdpb_inst_201_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2323 (
  .O(mux_o_2323),
  .I0(sdpb_inst_202_dout[18]),
  .I1(sdpb_inst_203_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2324 (
  .O(mux_o_2324),
  .I0(sdpb_inst_204_dout[18]),
  .I1(sdpb_inst_205_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2325 (
  .O(mux_o_2325),
  .I0(sdpb_inst_206_dout[18]),
  .I1(sdpb_inst_207_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2326 (
  .O(mux_o_2326),
  .I0(sdpb_inst_208_dout[18]),
  .I1(sdpb_inst_209_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2327 (
  .O(mux_o_2327),
  .I0(sdpb_inst_210_dout[18]),
  .I1(sdpb_inst_211_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2328 (
  .O(mux_o_2328),
  .I0(sdpb_inst_212_dout[18]),
  .I1(sdpb_inst_213_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2329 (
  .O(mux_o_2329),
  .I0(sdpb_inst_214_dout[18]),
  .I1(sdpb_inst_215_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2330 (
  .O(mux_o_2330),
  .I0(sdpb_inst_216_dout[18]),
  .I1(sdpb_inst_217_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2331 (
  .O(mux_o_2331),
  .I0(sdpb_inst_218_dout[18]),
  .I1(sdpb_inst_219_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2332 (
  .O(mux_o_2332),
  .I0(sdpb_inst_220_dout[18]),
  .I1(sdpb_inst_221_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2333 (
  .O(mux_o_2333),
  .I0(sdpb_inst_222_dout[18]),
  .I1(sdpb_inst_223_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2334 (
  .O(mux_o_2334),
  .I0(sdpb_inst_224_dout[18]),
  .I1(sdpb_inst_225_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2335 (
  .O(mux_o_2335),
  .I0(sdpb_inst_226_dout[18]),
  .I1(sdpb_inst_227_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2336 (
  .O(mux_o_2336),
  .I0(sdpb_inst_228_dout[18]),
  .I1(sdpb_inst_229_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2337 (
  .O(mux_o_2337),
  .I0(sdpb_inst_230_dout[18]),
  .I1(sdpb_inst_231_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2338 (
  .O(mux_o_2338),
  .I0(sdpb_inst_232_dout[18]),
  .I1(sdpb_inst_233_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2339 (
  .O(mux_o_2339),
  .I0(sdpb_inst_234_dout[18]),
  .I1(sdpb_inst_235_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2340 (
  .O(mux_o_2340),
  .I0(sdpb_inst_236_dout[18]),
  .I1(sdpb_inst_237_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2341 (
  .O(mux_o_2341),
  .I0(sdpb_inst_238_dout[18]),
  .I1(sdpb_inst_239_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2342 (
  .O(mux_o_2342),
  .I0(sdpb_inst_240_dout[18]),
  .I1(sdpb_inst_241_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2343 (
  .O(mux_o_2343),
  .I0(sdpb_inst_242_dout[18]),
  .I1(sdpb_inst_243_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2344 (
  .O(mux_o_2344),
  .I0(sdpb_inst_244_dout[18]),
  .I1(sdpb_inst_245_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2345 (
  .O(mux_o_2345),
  .I0(sdpb_inst_246_dout[18]),
  .I1(sdpb_inst_247_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2346 (
  .O(mux_o_2346),
  .I0(sdpb_inst_248_dout[18]),
  .I1(sdpb_inst_249_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2347 (
  .O(mux_o_2347),
  .I0(sdpb_inst_250_dout[18]),
  .I1(sdpb_inst_251_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2348 (
  .O(mux_o_2348),
  .I0(sdpb_inst_252_dout[18]),
  .I1(sdpb_inst_253_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2349 (
  .O(mux_o_2349),
  .I0(sdpb_inst_254_dout[18]),
  .I1(sdpb_inst_255_dout[18]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2350 (
  .O(mux_o_2350),
  .I0(mux_o_2286),
  .I1(mux_o_2287),
  .S0(dff_q_5)
);
MUX2 mux_inst_2351 (
  .O(mux_o_2351),
  .I0(mux_o_2288),
  .I1(mux_o_2289),
  .S0(dff_q_5)
);
MUX2 mux_inst_2352 (
  .O(mux_o_2352),
  .I0(mux_o_2290),
  .I1(mux_o_2291),
  .S0(dff_q_5)
);
MUX2 mux_inst_2353 (
  .O(mux_o_2353),
  .I0(mux_o_2292),
  .I1(mux_o_2293),
  .S0(dff_q_5)
);
MUX2 mux_inst_2354 (
  .O(mux_o_2354),
  .I0(mux_o_2294),
  .I1(mux_o_2295),
  .S0(dff_q_5)
);
MUX2 mux_inst_2355 (
  .O(mux_o_2355),
  .I0(mux_o_2296),
  .I1(mux_o_2297),
  .S0(dff_q_5)
);
MUX2 mux_inst_2356 (
  .O(mux_o_2356),
  .I0(mux_o_2298),
  .I1(mux_o_2299),
  .S0(dff_q_5)
);
MUX2 mux_inst_2357 (
  .O(mux_o_2357),
  .I0(mux_o_2300),
  .I1(mux_o_2301),
  .S0(dff_q_5)
);
MUX2 mux_inst_2358 (
  .O(mux_o_2358),
  .I0(mux_o_2302),
  .I1(mux_o_2303),
  .S0(dff_q_5)
);
MUX2 mux_inst_2359 (
  .O(mux_o_2359),
  .I0(mux_o_2304),
  .I1(mux_o_2305),
  .S0(dff_q_5)
);
MUX2 mux_inst_2360 (
  .O(mux_o_2360),
  .I0(mux_o_2306),
  .I1(mux_o_2307),
  .S0(dff_q_5)
);
MUX2 mux_inst_2361 (
  .O(mux_o_2361),
  .I0(mux_o_2308),
  .I1(mux_o_2309),
  .S0(dff_q_5)
);
MUX2 mux_inst_2362 (
  .O(mux_o_2362),
  .I0(mux_o_2310),
  .I1(mux_o_2311),
  .S0(dff_q_5)
);
MUX2 mux_inst_2363 (
  .O(mux_o_2363),
  .I0(mux_o_2312),
  .I1(mux_o_2313),
  .S0(dff_q_5)
);
MUX2 mux_inst_2364 (
  .O(mux_o_2364),
  .I0(mux_o_2314),
  .I1(mux_o_2315),
  .S0(dff_q_5)
);
MUX2 mux_inst_2365 (
  .O(mux_o_2365),
  .I0(mux_o_2316),
  .I1(mux_o_2317),
  .S0(dff_q_5)
);
MUX2 mux_inst_2366 (
  .O(mux_o_2366),
  .I0(mux_o_2318),
  .I1(mux_o_2319),
  .S0(dff_q_5)
);
MUX2 mux_inst_2367 (
  .O(mux_o_2367),
  .I0(mux_o_2320),
  .I1(mux_o_2321),
  .S0(dff_q_5)
);
MUX2 mux_inst_2368 (
  .O(mux_o_2368),
  .I0(mux_o_2322),
  .I1(mux_o_2323),
  .S0(dff_q_5)
);
MUX2 mux_inst_2369 (
  .O(mux_o_2369),
  .I0(mux_o_2324),
  .I1(mux_o_2325),
  .S0(dff_q_5)
);
MUX2 mux_inst_2370 (
  .O(mux_o_2370),
  .I0(mux_o_2326),
  .I1(mux_o_2327),
  .S0(dff_q_5)
);
MUX2 mux_inst_2371 (
  .O(mux_o_2371),
  .I0(mux_o_2328),
  .I1(mux_o_2329),
  .S0(dff_q_5)
);
MUX2 mux_inst_2372 (
  .O(mux_o_2372),
  .I0(mux_o_2330),
  .I1(mux_o_2331),
  .S0(dff_q_5)
);
MUX2 mux_inst_2373 (
  .O(mux_o_2373),
  .I0(mux_o_2332),
  .I1(mux_o_2333),
  .S0(dff_q_5)
);
MUX2 mux_inst_2374 (
  .O(mux_o_2374),
  .I0(mux_o_2334),
  .I1(mux_o_2335),
  .S0(dff_q_5)
);
MUX2 mux_inst_2375 (
  .O(mux_o_2375),
  .I0(mux_o_2336),
  .I1(mux_o_2337),
  .S0(dff_q_5)
);
MUX2 mux_inst_2376 (
  .O(mux_o_2376),
  .I0(mux_o_2338),
  .I1(mux_o_2339),
  .S0(dff_q_5)
);
MUX2 mux_inst_2377 (
  .O(mux_o_2377),
  .I0(mux_o_2340),
  .I1(mux_o_2341),
  .S0(dff_q_5)
);
MUX2 mux_inst_2378 (
  .O(mux_o_2378),
  .I0(mux_o_2342),
  .I1(mux_o_2343),
  .S0(dff_q_5)
);
MUX2 mux_inst_2379 (
  .O(mux_o_2379),
  .I0(mux_o_2344),
  .I1(mux_o_2345),
  .S0(dff_q_5)
);
MUX2 mux_inst_2380 (
  .O(mux_o_2380),
  .I0(mux_o_2346),
  .I1(mux_o_2347),
  .S0(dff_q_5)
);
MUX2 mux_inst_2381 (
  .O(mux_o_2381),
  .I0(mux_o_2348),
  .I1(mux_o_2349),
  .S0(dff_q_5)
);
MUX2 mux_inst_2382 (
  .O(mux_o_2382),
  .I0(mux_o_2350),
  .I1(mux_o_2351),
  .S0(dff_q_4)
);
MUX2 mux_inst_2383 (
  .O(mux_o_2383),
  .I0(mux_o_2352),
  .I1(mux_o_2353),
  .S0(dff_q_4)
);
MUX2 mux_inst_2384 (
  .O(mux_o_2384),
  .I0(mux_o_2354),
  .I1(mux_o_2355),
  .S0(dff_q_4)
);
MUX2 mux_inst_2385 (
  .O(mux_o_2385),
  .I0(mux_o_2356),
  .I1(mux_o_2357),
  .S0(dff_q_4)
);
MUX2 mux_inst_2386 (
  .O(mux_o_2386),
  .I0(mux_o_2358),
  .I1(mux_o_2359),
  .S0(dff_q_4)
);
MUX2 mux_inst_2387 (
  .O(mux_o_2387),
  .I0(mux_o_2360),
  .I1(mux_o_2361),
  .S0(dff_q_4)
);
MUX2 mux_inst_2388 (
  .O(mux_o_2388),
  .I0(mux_o_2362),
  .I1(mux_o_2363),
  .S0(dff_q_4)
);
MUX2 mux_inst_2389 (
  .O(mux_o_2389),
  .I0(mux_o_2364),
  .I1(mux_o_2365),
  .S0(dff_q_4)
);
MUX2 mux_inst_2390 (
  .O(mux_o_2390),
  .I0(mux_o_2366),
  .I1(mux_o_2367),
  .S0(dff_q_4)
);
MUX2 mux_inst_2391 (
  .O(mux_o_2391),
  .I0(mux_o_2368),
  .I1(mux_o_2369),
  .S0(dff_q_4)
);
MUX2 mux_inst_2392 (
  .O(mux_o_2392),
  .I0(mux_o_2370),
  .I1(mux_o_2371),
  .S0(dff_q_4)
);
MUX2 mux_inst_2393 (
  .O(mux_o_2393),
  .I0(mux_o_2372),
  .I1(mux_o_2373),
  .S0(dff_q_4)
);
MUX2 mux_inst_2394 (
  .O(mux_o_2394),
  .I0(mux_o_2374),
  .I1(mux_o_2375),
  .S0(dff_q_4)
);
MUX2 mux_inst_2395 (
  .O(mux_o_2395),
  .I0(mux_o_2376),
  .I1(mux_o_2377),
  .S0(dff_q_4)
);
MUX2 mux_inst_2396 (
  .O(mux_o_2396),
  .I0(mux_o_2378),
  .I1(mux_o_2379),
  .S0(dff_q_4)
);
MUX2 mux_inst_2397 (
  .O(mux_o_2397),
  .I0(mux_o_2380),
  .I1(mux_o_2381),
  .S0(dff_q_4)
);
MUX2 mux_inst_2398 (
  .O(mux_o_2398),
  .I0(mux_o_2382),
  .I1(mux_o_2383),
  .S0(dff_q_3)
);
MUX2 mux_inst_2399 (
  .O(mux_o_2399),
  .I0(mux_o_2384),
  .I1(mux_o_2385),
  .S0(dff_q_3)
);
MUX2 mux_inst_2400 (
  .O(mux_o_2400),
  .I0(mux_o_2386),
  .I1(mux_o_2387),
  .S0(dff_q_3)
);
MUX2 mux_inst_2401 (
  .O(mux_o_2401),
  .I0(mux_o_2388),
  .I1(mux_o_2389),
  .S0(dff_q_3)
);
MUX2 mux_inst_2402 (
  .O(mux_o_2402),
  .I0(mux_o_2390),
  .I1(mux_o_2391),
  .S0(dff_q_3)
);
MUX2 mux_inst_2403 (
  .O(mux_o_2403),
  .I0(mux_o_2392),
  .I1(mux_o_2393),
  .S0(dff_q_3)
);
MUX2 mux_inst_2404 (
  .O(mux_o_2404),
  .I0(mux_o_2394),
  .I1(mux_o_2395),
  .S0(dff_q_3)
);
MUX2 mux_inst_2405 (
  .O(mux_o_2405),
  .I0(mux_o_2396),
  .I1(mux_o_2397),
  .S0(dff_q_3)
);
MUX2 mux_inst_2406 (
  .O(mux_o_2406),
  .I0(mux_o_2398),
  .I1(mux_o_2399),
  .S0(dff_q_2)
);
MUX2 mux_inst_2407 (
  .O(mux_o_2407),
  .I0(mux_o_2400),
  .I1(mux_o_2401),
  .S0(dff_q_2)
);
MUX2 mux_inst_2408 (
  .O(mux_o_2408),
  .I0(mux_o_2402),
  .I1(mux_o_2403),
  .S0(dff_q_2)
);
MUX2 mux_inst_2409 (
  .O(mux_o_2409),
  .I0(mux_o_2404),
  .I1(mux_o_2405),
  .S0(dff_q_2)
);
MUX2 mux_inst_2410 (
  .O(mux_o_2410),
  .I0(mux_o_2406),
  .I1(mux_o_2407),
  .S0(dff_q_1)
);
MUX2 mux_inst_2411 (
  .O(mux_o_2411),
  .I0(mux_o_2408),
  .I1(mux_o_2409),
  .S0(dff_q_1)
);
MUX2 mux_inst_2412 (
  .O(dout[18]),
  .I0(mux_o_2410),
  .I1(mux_o_2411),
  .S0(dff_q_0)
);
MUX2 mux_inst_2413 (
  .O(mux_o_2413),
  .I0(sdpb_inst_128_dout[19]),
  .I1(sdpb_inst_129_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2414 (
  .O(mux_o_2414),
  .I0(sdpb_inst_130_dout[19]),
  .I1(sdpb_inst_131_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2415 (
  .O(mux_o_2415),
  .I0(sdpb_inst_132_dout[19]),
  .I1(sdpb_inst_133_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2416 (
  .O(mux_o_2416),
  .I0(sdpb_inst_134_dout[19]),
  .I1(sdpb_inst_135_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2417 (
  .O(mux_o_2417),
  .I0(sdpb_inst_136_dout[19]),
  .I1(sdpb_inst_137_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2418 (
  .O(mux_o_2418),
  .I0(sdpb_inst_138_dout[19]),
  .I1(sdpb_inst_139_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2419 (
  .O(mux_o_2419),
  .I0(sdpb_inst_140_dout[19]),
  .I1(sdpb_inst_141_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2420 (
  .O(mux_o_2420),
  .I0(sdpb_inst_142_dout[19]),
  .I1(sdpb_inst_143_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2421 (
  .O(mux_o_2421),
  .I0(sdpb_inst_144_dout[19]),
  .I1(sdpb_inst_145_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2422 (
  .O(mux_o_2422),
  .I0(sdpb_inst_146_dout[19]),
  .I1(sdpb_inst_147_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2423 (
  .O(mux_o_2423),
  .I0(sdpb_inst_148_dout[19]),
  .I1(sdpb_inst_149_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2424 (
  .O(mux_o_2424),
  .I0(sdpb_inst_150_dout[19]),
  .I1(sdpb_inst_151_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2425 (
  .O(mux_o_2425),
  .I0(sdpb_inst_152_dout[19]),
  .I1(sdpb_inst_153_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2426 (
  .O(mux_o_2426),
  .I0(sdpb_inst_154_dout[19]),
  .I1(sdpb_inst_155_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2427 (
  .O(mux_o_2427),
  .I0(sdpb_inst_156_dout[19]),
  .I1(sdpb_inst_157_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2428 (
  .O(mux_o_2428),
  .I0(sdpb_inst_158_dout[19]),
  .I1(sdpb_inst_159_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2429 (
  .O(mux_o_2429),
  .I0(sdpb_inst_160_dout[19]),
  .I1(sdpb_inst_161_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2430 (
  .O(mux_o_2430),
  .I0(sdpb_inst_162_dout[19]),
  .I1(sdpb_inst_163_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2431 (
  .O(mux_o_2431),
  .I0(sdpb_inst_164_dout[19]),
  .I1(sdpb_inst_165_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2432 (
  .O(mux_o_2432),
  .I0(sdpb_inst_166_dout[19]),
  .I1(sdpb_inst_167_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2433 (
  .O(mux_o_2433),
  .I0(sdpb_inst_168_dout[19]),
  .I1(sdpb_inst_169_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2434 (
  .O(mux_o_2434),
  .I0(sdpb_inst_170_dout[19]),
  .I1(sdpb_inst_171_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2435 (
  .O(mux_o_2435),
  .I0(sdpb_inst_172_dout[19]),
  .I1(sdpb_inst_173_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2436 (
  .O(mux_o_2436),
  .I0(sdpb_inst_174_dout[19]),
  .I1(sdpb_inst_175_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2437 (
  .O(mux_o_2437),
  .I0(sdpb_inst_176_dout[19]),
  .I1(sdpb_inst_177_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2438 (
  .O(mux_o_2438),
  .I0(sdpb_inst_178_dout[19]),
  .I1(sdpb_inst_179_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2439 (
  .O(mux_o_2439),
  .I0(sdpb_inst_180_dout[19]),
  .I1(sdpb_inst_181_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2440 (
  .O(mux_o_2440),
  .I0(sdpb_inst_182_dout[19]),
  .I1(sdpb_inst_183_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2441 (
  .O(mux_o_2441),
  .I0(sdpb_inst_184_dout[19]),
  .I1(sdpb_inst_185_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2442 (
  .O(mux_o_2442),
  .I0(sdpb_inst_186_dout[19]),
  .I1(sdpb_inst_187_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2443 (
  .O(mux_o_2443),
  .I0(sdpb_inst_188_dout[19]),
  .I1(sdpb_inst_189_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2444 (
  .O(mux_o_2444),
  .I0(sdpb_inst_190_dout[19]),
  .I1(sdpb_inst_191_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2445 (
  .O(mux_o_2445),
  .I0(sdpb_inst_192_dout[19]),
  .I1(sdpb_inst_193_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2446 (
  .O(mux_o_2446),
  .I0(sdpb_inst_194_dout[19]),
  .I1(sdpb_inst_195_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2447 (
  .O(mux_o_2447),
  .I0(sdpb_inst_196_dout[19]),
  .I1(sdpb_inst_197_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2448 (
  .O(mux_o_2448),
  .I0(sdpb_inst_198_dout[19]),
  .I1(sdpb_inst_199_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2449 (
  .O(mux_o_2449),
  .I0(sdpb_inst_200_dout[19]),
  .I1(sdpb_inst_201_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2450 (
  .O(mux_o_2450),
  .I0(sdpb_inst_202_dout[19]),
  .I1(sdpb_inst_203_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2451 (
  .O(mux_o_2451),
  .I0(sdpb_inst_204_dout[19]),
  .I1(sdpb_inst_205_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2452 (
  .O(mux_o_2452),
  .I0(sdpb_inst_206_dout[19]),
  .I1(sdpb_inst_207_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2453 (
  .O(mux_o_2453),
  .I0(sdpb_inst_208_dout[19]),
  .I1(sdpb_inst_209_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2454 (
  .O(mux_o_2454),
  .I0(sdpb_inst_210_dout[19]),
  .I1(sdpb_inst_211_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2455 (
  .O(mux_o_2455),
  .I0(sdpb_inst_212_dout[19]),
  .I1(sdpb_inst_213_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2456 (
  .O(mux_o_2456),
  .I0(sdpb_inst_214_dout[19]),
  .I1(sdpb_inst_215_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2457 (
  .O(mux_o_2457),
  .I0(sdpb_inst_216_dout[19]),
  .I1(sdpb_inst_217_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2458 (
  .O(mux_o_2458),
  .I0(sdpb_inst_218_dout[19]),
  .I1(sdpb_inst_219_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2459 (
  .O(mux_o_2459),
  .I0(sdpb_inst_220_dout[19]),
  .I1(sdpb_inst_221_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2460 (
  .O(mux_o_2460),
  .I0(sdpb_inst_222_dout[19]),
  .I1(sdpb_inst_223_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2461 (
  .O(mux_o_2461),
  .I0(sdpb_inst_224_dout[19]),
  .I1(sdpb_inst_225_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2462 (
  .O(mux_o_2462),
  .I0(sdpb_inst_226_dout[19]),
  .I1(sdpb_inst_227_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2463 (
  .O(mux_o_2463),
  .I0(sdpb_inst_228_dout[19]),
  .I1(sdpb_inst_229_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2464 (
  .O(mux_o_2464),
  .I0(sdpb_inst_230_dout[19]),
  .I1(sdpb_inst_231_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2465 (
  .O(mux_o_2465),
  .I0(sdpb_inst_232_dout[19]),
  .I1(sdpb_inst_233_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2466 (
  .O(mux_o_2466),
  .I0(sdpb_inst_234_dout[19]),
  .I1(sdpb_inst_235_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2467 (
  .O(mux_o_2467),
  .I0(sdpb_inst_236_dout[19]),
  .I1(sdpb_inst_237_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2468 (
  .O(mux_o_2468),
  .I0(sdpb_inst_238_dout[19]),
  .I1(sdpb_inst_239_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2469 (
  .O(mux_o_2469),
  .I0(sdpb_inst_240_dout[19]),
  .I1(sdpb_inst_241_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2470 (
  .O(mux_o_2470),
  .I0(sdpb_inst_242_dout[19]),
  .I1(sdpb_inst_243_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2471 (
  .O(mux_o_2471),
  .I0(sdpb_inst_244_dout[19]),
  .I1(sdpb_inst_245_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2472 (
  .O(mux_o_2472),
  .I0(sdpb_inst_246_dout[19]),
  .I1(sdpb_inst_247_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2473 (
  .O(mux_o_2473),
  .I0(sdpb_inst_248_dout[19]),
  .I1(sdpb_inst_249_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2474 (
  .O(mux_o_2474),
  .I0(sdpb_inst_250_dout[19]),
  .I1(sdpb_inst_251_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2475 (
  .O(mux_o_2475),
  .I0(sdpb_inst_252_dout[19]),
  .I1(sdpb_inst_253_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2476 (
  .O(mux_o_2476),
  .I0(sdpb_inst_254_dout[19]),
  .I1(sdpb_inst_255_dout[19]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2477 (
  .O(mux_o_2477),
  .I0(mux_o_2413),
  .I1(mux_o_2414),
  .S0(dff_q_5)
);
MUX2 mux_inst_2478 (
  .O(mux_o_2478),
  .I0(mux_o_2415),
  .I1(mux_o_2416),
  .S0(dff_q_5)
);
MUX2 mux_inst_2479 (
  .O(mux_o_2479),
  .I0(mux_o_2417),
  .I1(mux_o_2418),
  .S0(dff_q_5)
);
MUX2 mux_inst_2480 (
  .O(mux_o_2480),
  .I0(mux_o_2419),
  .I1(mux_o_2420),
  .S0(dff_q_5)
);
MUX2 mux_inst_2481 (
  .O(mux_o_2481),
  .I0(mux_o_2421),
  .I1(mux_o_2422),
  .S0(dff_q_5)
);
MUX2 mux_inst_2482 (
  .O(mux_o_2482),
  .I0(mux_o_2423),
  .I1(mux_o_2424),
  .S0(dff_q_5)
);
MUX2 mux_inst_2483 (
  .O(mux_o_2483),
  .I0(mux_o_2425),
  .I1(mux_o_2426),
  .S0(dff_q_5)
);
MUX2 mux_inst_2484 (
  .O(mux_o_2484),
  .I0(mux_o_2427),
  .I1(mux_o_2428),
  .S0(dff_q_5)
);
MUX2 mux_inst_2485 (
  .O(mux_o_2485),
  .I0(mux_o_2429),
  .I1(mux_o_2430),
  .S0(dff_q_5)
);
MUX2 mux_inst_2486 (
  .O(mux_o_2486),
  .I0(mux_o_2431),
  .I1(mux_o_2432),
  .S0(dff_q_5)
);
MUX2 mux_inst_2487 (
  .O(mux_o_2487),
  .I0(mux_o_2433),
  .I1(mux_o_2434),
  .S0(dff_q_5)
);
MUX2 mux_inst_2488 (
  .O(mux_o_2488),
  .I0(mux_o_2435),
  .I1(mux_o_2436),
  .S0(dff_q_5)
);
MUX2 mux_inst_2489 (
  .O(mux_o_2489),
  .I0(mux_o_2437),
  .I1(mux_o_2438),
  .S0(dff_q_5)
);
MUX2 mux_inst_2490 (
  .O(mux_o_2490),
  .I0(mux_o_2439),
  .I1(mux_o_2440),
  .S0(dff_q_5)
);
MUX2 mux_inst_2491 (
  .O(mux_o_2491),
  .I0(mux_o_2441),
  .I1(mux_o_2442),
  .S0(dff_q_5)
);
MUX2 mux_inst_2492 (
  .O(mux_o_2492),
  .I0(mux_o_2443),
  .I1(mux_o_2444),
  .S0(dff_q_5)
);
MUX2 mux_inst_2493 (
  .O(mux_o_2493),
  .I0(mux_o_2445),
  .I1(mux_o_2446),
  .S0(dff_q_5)
);
MUX2 mux_inst_2494 (
  .O(mux_o_2494),
  .I0(mux_o_2447),
  .I1(mux_o_2448),
  .S0(dff_q_5)
);
MUX2 mux_inst_2495 (
  .O(mux_o_2495),
  .I0(mux_o_2449),
  .I1(mux_o_2450),
  .S0(dff_q_5)
);
MUX2 mux_inst_2496 (
  .O(mux_o_2496),
  .I0(mux_o_2451),
  .I1(mux_o_2452),
  .S0(dff_q_5)
);
MUX2 mux_inst_2497 (
  .O(mux_o_2497),
  .I0(mux_o_2453),
  .I1(mux_o_2454),
  .S0(dff_q_5)
);
MUX2 mux_inst_2498 (
  .O(mux_o_2498),
  .I0(mux_o_2455),
  .I1(mux_o_2456),
  .S0(dff_q_5)
);
MUX2 mux_inst_2499 (
  .O(mux_o_2499),
  .I0(mux_o_2457),
  .I1(mux_o_2458),
  .S0(dff_q_5)
);
MUX2 mux_inst_2500 (
  .O(mux_o_2500),
  .I0(mux_o_2459),
  .I1(mux_o_2460),
  .S0(dff_q_5)
);
MUX2 mux_inst_2501 (
  .O(mux_o_2501),
  .I0(mux_o_2461),
  .I1(mux_o_2462),
  .S0(dff_q_5)
);
MUX2 mux_inst_2502 (
  .O(mux_o_2502),
  .I0(mux_o_2463),
  .I1(mux_o_2464),
  .S0(dff_q_5)
);
MUX2 mux_inst_2503 (
  .O(mux_o_2503),
  .I0(mux_o_2465),
  .I1(mux_o_2466),
  .S0(dff_q_5)
);
MUX2 mux_inst_2504 (
  .O(mux_o_2504),
  .I0(mux_o_2467),
  .I1(mux_o_2468),
  .S0(dff_q_5)
);
MUX2 mux_inst_2505 (
  .O(mux_o_2505),
  .I0(mux_o_2469),
  .I1(mux_o_2470),
  .S0(dff_q_5)
);
MUX2 mux_inst_2506 (
  .O(mux_o_2506),
  .I0(mux_o_2471),
  .I1(mux_o_2472),
  .S0(dff_q_5)
);
MUX2 mux_inst_2507 (
  .O(mux_o_2507),
  .I0(mux_o_2473),
  .I1(mux_o_2474),
  .S0(dff_q_5)
);
MUX2 mux_inst_2508 (
  .O(mux_o_2508),
  .I0(mux_o_2475),
  .I1(mux_o_2476),
  .S0(dff_q_5)
);
MUX2 mux_inst_2509 (
  .O(mux_o_2509),
  .I0(mux_o_2477),
  .I1(mux_o_2478),
  .S0(dff_q_4)
);
MUX2 mux_inst_2510 (
  .O(mux_o_2510),
  .I0(mux_o_2479),
  .I1(mux_o_2480),
  .S0(dff_q_4)
);
MUX2 mux_inst_2511 (
  .O(mux_o_2511),
  .I0(mux_o_2481),
  .I1(mux_o_2482),
  .S0(dff_q_4)
);
MUX2 mux_inst_2512 (
  .O(mux_o_2512),
  .I0(mux_o_2483),
  .I1(mux_o_2484),
  .S0(dff_q_4)
);
MUX2 mux_inst_2513 (
  .O(mux_o_2513),
  .I0(mux_o_2485),
  .I1(mux_o_2486),
  .S0(dff_q_4)
);
MUX2 mux_inst_2514 (
  .O(mux_o_2514),
  .I0(mux_o_2487),
  .I1(mux_o_2488),
  .S0(dff_q_4)
);
MUX2 mux_inst_2515 (
  .O(mux_o_2515),
  .I0(mux_o_2489),
  .I1(mux_o_2490),
  .S0(dff_q_4)
);
MUX2 mux_inst_2516 (
  .O(mux_o_2516),
  .I0(mux_o_2491),
  .I1(mux_o_2492),
  .S0(dff_q_4)
);
MUX2 mux_inst_2517 (
  .O(mux_o_2517),
  .I0(mux_o_2493),
  .I1(mux_o_2494),
  .S0(dff_q_4)
);
MUX2 mux_inst_2518 (
  .O(mux_o_2518),
  .I0(mux_o_2495),
  .I1(mux_o_2496),
  .S0(dff_q_4)
);
MUX2 mux_inst_2519 (
  .O(mux_o_2519),
  .I0(mux_o_2497),
  .I1(mux_o_2498),
  .S0(dff_q_4)
);
MUX2 mux_inst_2520 (
  .O(mux_o_2520),
  .I0(mux_o_2499),
  .I1(mux_o_2500),
  .S0(dff_q_4)
);
MUX2 mux_inst_2521 (
  .O(mux_o_2521),
  .I0(mux_o_2501),
  .I1(mux_o_2502),
  .S0(dff_q_4)
);
MUX2 mux_inst_2522 (
  .O(mux_o_2522),
  .I0(mux_o_2503),
  .I1(mux_o_2504),
  .S0(dff_q_4)
);
MUX2 mux_inst_2523 (
  .O(mux_o_2523),
  .I0(mux_o_2505),
  .I1(mux_o_2506),
  .S0(dff_q_4)
);
MUX2 mux_inst_2524 (
  .O(mux_o_2524),
  .I0(mux_o_2507),
  .I1(mux_o_2508),
  .S0(dff_q_4)
);
MUX2 mux_inst_2525 (
  .O(mux_o_2525),
  .I0(mux_o_2509),
  .I1(mux_o_2510),
  .S0(dff_q_3)
);
MUX2 mux_inst_2526 (
  .O(mux_o_2526),
  .I0(mux_o_2511),
  .I1(mux_o_2512),
  .S0(dff_q_3)
);
MUX2 mux_inst_2527 (
  .O(mux_o_2527),
  .I0(mux_o_2513),
  .I1(mux_o_2514),
  .S0(dff_q_3)
);
MUX2 mux_inst_2528 (
  .O(mux_o_2528),
  .I0(mux_o_2515),
  .I1(mux_o_2516),
  .S0(dff_q_3)
);
MUX2 mux_inst_2529 (
  .O(mux_o_2529),
  .I0(mux_o_2517),
  .I1(mux_o_2518),
  .S0(dff_q_3)
);
MUX2 mux_inst_2530 (
  .O(mux_o_2530),
  .I0(mux_o_2519),
  .I1(mux_o_2520),
  .S0(dff_q_3)
);
MUX2 mux_inst_2531 (
  .O(mux_o_2531),
  .I0(mux_o_2521),
  .I1(mux_o_2522),
  .S0(dff_q_3)
);
MUX2 mux_inst_2532 (
  .O(mux_o_2532),
  .I0(mux_o_2523),
  .I1(mux_o_2524),
  .S0(dff_q_3)
);
MUX2 mux_inst_2533 (
  .O(mux_o_2533),
  .I0(mux_o_2525),
  .I1(mux_o_2526),
  .S0(dff_q_2)
);
MUX2 mux_inst_2534 (
  .O(mux_o_2534),
  .I0(mux_o_2527),
  .I1(mux_o_2528),
  .S0(dff_q_2)
);
MUX2 mux_inst_2535 (
  .O(mux_o_2535),
  .I0(mux_o_2529),
  .I1(mux_o_2530),
  .S0(dff_q_2)
);
MUX2 mux_inst_2536 (
  .O(mux_o_2536),
  .I0(mux_o_2531),
  .I1(mux_o_2532),
  .S0(dff_q_2)
);
MUX2 mux_inst_2537 (
  .O(mux_o_2537),
  .I0(mux_o_2533),
  .I1(mux_o_2534),
  .S0(dff_q_1)
);
MUX2 mux_inst_2538 (
  .O(mux_o_2538),
  .I0(mux_o_2535),
  .I1(mux_o_2536),
  .S0(dff_q_1)
);
MUX2 mux_inst_2539 (
  .O(dout[19]),
  .I0(mux_o_2537),
  .I1(mux_o_2538),
  .S0(dff_q_0)
);
MUX2 mux_inst_2540 (
  .O(mux_o_2540),
  .I0(sdpb_inst_128_dout[20]),
  .I1(sdpb_inst_129_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2541 (
  .O(mux_o_2541),
  .I0(sdpb_inst_130_dout[20]),
  .I1(sdpb_inst_131_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2542 (
  .O(mux_o_2542),
  .I0(sdpb_inst_132_dout[20]),
  .I1(sdpb_inst_133_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2543 (
  .O(mux_o_2543),
  .I0(sdpb_inst_134_dout[20]),
  .I1(sdpb_inst_135_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2544 (
  .O(mux_o_2544),
  .I0(sdpb_inst_136_dout[20]),
  .I1(sdpb_inst_137_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2545 (
  .O(mux_o_2545),
  .I0(sdpb_inst_138_dout[20]),
  .I1(sdpb_inst_139_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2546 (
  .O(mux_o_2546),
  .I0(sdpb_inst_140_dout[20]),
  .I1(sdpb_inst_141_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2547 (
  .O(mux_o_2547),
  .I0(sdpb_inst_142_dout[20]),
  .I1(sdpb_inst_143_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2548 (
  .O(mux_o_2548),
  .I0(sdpb_inst_144_dout[20]),
  .I1(sdpb_inst_145_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2549 (
  .O(mux_o_2549),
  .I0(sdpb_inst_146_dout[20]),
  .I1(sdpb_inst_147_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2550 (
  .O(mux_o_2550),
  .I0(sdpb_inst_148_dout[20]),
  .I1(sdpb_inst_149_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2551 (
  .O(mux_o_2551),
  .I0(sdpb_inst_150_dout[20]),
  .I1(sdpb_inst_151_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2552 (
  .O(mux_o_2552),
  .I0(sdpb_inst_152_dout[20]),
  .I1(sdpb_inst_153_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2553 (
  .O(mux_o_2553),
  .I0(sdpb_inst_154_dout[20]),
  .I1(sdpb_inst_155_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2554 (
  .O(mux_o_2554),
  .I0(sdpb_inst_156_dout[20]),
  .I1(sdpb_inst_157_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2555 (
  .O(mux_o_2555),
  .I0(sdpb_inst_158_dout[20]),
  .I1(sdpb_inst_159_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2556 (
  .O(mux_o_2556),
  .I0(sdpb_inst_160_dout[20]),
  .I1(sdpb_inst_161_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2557 (
  .O(mux_o_2557),
  .I0(sdpb_inst_162_dout[20]),
  .I1(sdpb_inst_163_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2558 (
  .O(mux_o_2558),
  .I0(sdpb_inst_164_dout[20]),
  .I1(sdpb_inst_165_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2559 (
  .O(mux_o_2559),
  .I0(sdpb_inst_166_dout[20]),
  .I1(sdpb_inst_167_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2560 (
  .O(mux_o_2560),
  .I0(sdpb_inst_168_dout[20]),
  .I1(sdpb_inst_169_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2561 (
  .O(mux_o_2561),
  .I0(sdpb_inst_170_dout[20]),
  .I1(sdpb_inst_171_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2562 (
  .O(mux_o_2562),
  .I0(sdpb_inst_172_dout[20]),
  .I1(sdpb_inst_173_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2563 (
  .O(mux_o_2563),
  .I0(sdpb_inst_174_dout[20]),
  .I1(sdpb_inst_175_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2564 (
  .O(mux_o_2564),
  .I0(sdpb_inst_176_dout[20]),
  .I1(sdpb_inst_177_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2565 (
  .O(mux_o_2565),
  .I0(sdpb_inst_178_dout[20]),
  .I1(sdpb_inst_179_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2566 (
  .O(mux_o_2566),
  .I0(sdpb_inst_180_dout[20]),
  .I1(sdpb_inst_181_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2567 (
  .O(mux_o_2567),
  .I0(sdpb_inst_182_dout[20]),
  .I1(sdpb_inst_183_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2568 (
  .O(mux_o_2568),
  .I0(sdpb_inst_184_dout[20]),
  .I1(sdpb_inst_185_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2569 (
  .O(mux_o_2569),
  .I0(sdpb_inst_186_dout[20]),
  .I1(sdpb_inst_187_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2570 (
  .O(mux_o_2570),
  .I0(sdpb_inst_188_dout[20]),
  .I1(sdpb_inst_189_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2571 (
  .O(mux_o_2571),
  .I0(sdpb_inst_190_dout[20]),
  .I1(sdpb_inst_191_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2572 (
  .O(mux_o_2572),
  .I0(sdpb_inst_192_dout[20]),
  .I1(sdpb_inst_193_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2573 (
  .O(mux_o_2573),
  .I0(sdpb_inst_194_dout[20]),
  .I1(sdpb_inst_195_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2574 (
  .O(mux_o_2574),
  .I0(sdpb_inst_196_dout[20]),
  .I1(sdpb_inst_197_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2575 (
  .O(mux_o_2575),
  .I0(sdpb_inst_198_dout[20]),
  .I1(sdpb_inst_199_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2576 (
  .O(mux_o_2576),
  .I0(sdpb_inst_200_dout[20]),
  .I1(sdpb_inst_201_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2577 (
  .O(mux_o_2577),
  .I0(sdpb_inst_202_dout[20]),
  .I1(sdpb_inst_203_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2578 (
  .O(mux_o_2578),
  .I0(sdpb_inst_204_dout[20]),
  .I1(sdpb_inst_205_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2579 (
  .O(mux_o_2579),
  .I0(sdpb_inst_206_dout[20]),
  .I1(sdpb_inst_207_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2580 (
  .O(mux_o_2580),
  .I0(sdpb_inst_208_dout[20]),
  .I1(sdpb_inst_209_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2581 (
  .O(mux_o_2581),
  .I0(sdpb_inst_210_dout[20]),
  .I1(sdpb_inst_211_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2582 (
  .O(mux_o_2582),
  .I0(sdpb_inst_212_dout[20]),
  .I1(sdpb_inst_213_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2583 (
  .O(mux_o_2583),
  .I0(sdpb_inst_214_dout[20]),
  .I1(sdpb_inst_215_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2584 (
  .O(mux_o_2584),
  .I0(sdpb_inst_216_dout[20]),
  .I1(sdpb_inst_217_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2585 (
  .O(mux_o_2585),
  .I0(sdpb_inst_218_dout[20]),
  .I1(sdpb_inst_219_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2586 (
  .O(mux_o_2586),
  .I0(sdpb_inst_220_dout[20]),
  .I1(sdpb_inst_221_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2587 (
  .O(mux_o_2587),
  .I0(sdpb_inst_222_dout[20]),
  .I1(sdpb_inst_223_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2588 (
  .O(mux_o_2588),
  .I0(sdpb_inst_224_dout[20]),
  .I1(sdpb_inst_225_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2589 (
  .O(mux_o_2589),
  .I0(sdpb_inst_226_dout[20]),
  .I1(sdpb_inst_227_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2590 (
  .O(mux_o_2590),
  .I0(sdpb_inst_228_dout[20]),
  .I1(sdpb_inst_229_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2591 (
  .O(mux_o_2591),
  .I0(sdpb_inst_230_dout[20]),
  .I1(sdpb_inst_231_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2592 (
  .O(mux_o_2592),
  .I0(sdpb_inst_232_dout[20]),
  .I1(sdpb_inst_233_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2593 (
  .O(mux_o_2593),
  .I0(sdpb_inst_234_dout[20]),
  .I1(sdpb_inst_235_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2594 (
  .O(mux_o_2594),
  .I0(sdpb_inst_236_dout[20]),
  .I1(sdpb_inst_237_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2595 (
  .O(mux_o_2595),
  .I0(sdpb_inst_238_dout[20]),
  .I1(sdpb_inst_239_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2596 (
  .O(mux_o_2596),
  .I0(sdpb_inst_240_dout[20]),
  .I1(sdpb_inst_241_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2597 (
  .O(mux_o_2597),
  .I0(sdpb_inst_242_dout[20]),
  .I1(sdpb_inst_243_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2598 (
  .O(mux_o_2598),
  .I0(sdpb_inst_244_dout[20]),
  .I1(sdpb_inst_245_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2599 (
  .O(mux_o_2599),
  .I0(sdpb_inst_246_dout[20]),
  .I1(sdpb_inst_247_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2600 (
  .O(mux_o_2600),
  .I0(sdpb_inst_248_dout[20]),
  .I1(sdpb_inst_249_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2601 (
  .O(mux_o_2601),
  .I0(sdpb_inst_250_dout[20]),
  .I1(sdpb_inst_251_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2602 (
  .O(mux_o_2602),
  .I0(sdpb_inst_252_dout[20]),
  .I1(sdpb_inst_253_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2603 (
  .O(mux_o_2603),
  .I0(sdpb_inst_254_dout[20]),
  .I1(sdpb_inst_255_dout[20]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2604 (
  .O(mux_o_2604),
  .I0(mux_o_2540),
  .I1(mux_o_2541),
  .S0(dff_q_5)
);
MUX2 mux_inst_2605 (
  .O(mux_o_2605),
  .I0(mux_o_2542),
  .I1(mux_o_2543),
  .S0(dff_q_5)
);
MUX2 mux_inst_2606 (
  .O(mux_o_2606),
  .I0(mux_o_2544),
  .I1(mux_o_2545),
  .S0(dff_q_5)
);
MUX2 mux_inst_2607 (
  .O(mux_o_2607),
  .I0(mux_o_2546),
  .I1(mux_o_2547),
  .S0(dff_q_5)
);
MUX2 mux_inst_2608 (
  .O(mux_o_2608),
  .I0(mux_o_2548),
  .I1(mux_o_2549),
  .S0(dff_q_5)
);
MUX2 mux_inst_2609 (
  .O(mux_o_2609),
  .I0(mux_o_2550),
  .I1(mux_o_2551),
  .S0(dff_q_5)
);
MUX2 mux_inst_2610 (
  .O(mux_o_2610),
  .I0(mux_o_2552),
  .I1(mux_o_2553),
  .S0(dff_q_5)
);
MUX2 mux_inst_2611 (
  .O(mux_o_2611),
  .I0(mux_o_2554),
  .I1(mux_o_2555),
  .S0(dff_q_5)
);
MUX2 mux_inst_2612 (
  .O(mux_o_2612),
  .I0(mux_o_2556),
  .I1(mux_o_2557),
  .S0(dff_q_5)
);
MUX2 mux_inst_2613 (
  .O(mux_o_2613),
  .I0(mux_o_2558),
  .I1(mux_o_2559),
  .S0(dff_q_5)
);
MUX2 mux_inst_2614 (
  .O(mux_o_2614),
  .I0(mux_o_2560),
  .I1(mux_o_2561),
  .S0(dff_q_5)
);
MUX2 mux_inst_2615 (
  .O(mux_o_2615),
  .I0(mux_o_2562),
  .I1(mux_o_2563),
  .S0(dff_q_5)
);
MUX2 mux_inst_2616 (
  .O(mux_o_2616),
  .I0(mux_o_2564),
  .I1(mux_o_2565),
  .S0(dff_q_5)
);
MUX2 mux_inst_2617 (
  .O(mux_o_2617),
  .I0(mux_o_2566),
  .I1(mux_o_2567),
  .S0(dff_q_5)
);
MUX2 mux_inst_2618 (
  .O(mux_o_2618),
  .I0(mux_o_2568),
  .I1(mux_o_2569),
  .S0(dff_q_5)
);
MUX2 mux_inst_2619 (
  .O(mux_o_2619),
  .I0(mux_o_2570),
  .I1(mux_o_2571),
  .S0(dff_q_5)
);
MUX2 mux_inst_2620 (
  .O(mux_o_2620),
  .I0(mux_o_2572),
  .I1(mux_o_2573),
  .S0(dff_q_5)
);
MUX2 mux_inst_2621 (
  .O(mux_o_2621),
  .I0(mux_o_2574),
  .I1(mux_o_2575),
  .S0(dff_q_5)
);
MUX2 mux_inst_2622 (
  .O(mux_o_2622),
  .I0(mux_o_2576),
  .I1(mux_o_2577),
  .S0(dff_q_5)
);
MUX2 mux_inst_2623 (
  .O(mux_o_2623),
  .I0(mux_o_2578),
  .I1(mux_o_2579),
  .S0(dff_q_5)
);
MUX2 mux_inst_2624 (
  .O(mux_o_2624),
  .I0(mux_o_2580),
  .I1(mux_o_2581),
  .S0(dff_q_5)
);
MUX2 mux_inst_2625 (
  .O(mux_o_2625),
  .I0(mux_o_2582),
  .I1(mux_o_2583),
  .S0(dff_q_5)
);
MUX2 mux_inst_2626 (
  .O(mux_o_2626),
  .I0(mux_o_2584),
  .I1(mux_o_2585),
  .S0(dff_q_5)
);
MUX2 mux_inst_2627 (
  .O(mux_o_2627),
  .I0(mux_o_2586),
  .I1(mux_o_2587),
  .S0(dff_q_5)
);
MUX2 mux_inst_2628 (
  .O(mux_o_2628),
  .I0(mux_o_2588),
  .I1(mux_o_2589),
  .S0(dff_q_5)
);
MUX2 mux_inst_2629 (
  .O(mux_o_2629),
  .I0(mux_o_2590),
  .I1(mux_o_2591),
  .S0(dff_q_5)
);
MUX2 mux_inst_2630 (
  .O(mux_o_2630),
  .I0(mux_o_2592),
  .I1(mux_o_2593),
  .S0(dff_q_5)
);
MUX2 mux_inst_2631 (
  .O(mux_o_2631),
  .I0(mux_o_2594),
  .I1(mux_o_2595),
  .S0(dff_q_5)
);
MUX2 mux_inst_2632 (
  .O(mux_o_2632),
  .I0(mux_o_2596),
  .I1(mux_o_2597),
  .S0(dff_q_5)
);
MUX2 mux_inst_2633 (
  .O(mux_o_2633),
  .I0(mux_o_2598),
  .I1(mux_o_2599),
  .S0(dff_q_5)
);
MUX2 mux_inst_2634 (
  .O(mux_o_2634),
  .I0(mux_o_2600),
  .I1(mux_o_2601),
  .S0(dff_q_5)
);
MUX2 mux_inst_2635 (
  .O(mux_o_2635),
  .I0(mux_o_2602),
  .I1(mux_o_2603),
  .S0(dff_q_5)
);
MUX2 mux_inst_2636 (
  .O(mux_o_2636),
  .I0(mux_o_2604),
  .I1(mux_o_2605),
  .S0(dff_q_4)
);
MUX2 mux_inst_2637 (
  .O(mux_o_2637),
  .I0(mux_o_2606),
  .I1(mux_o_2607),
  .S0(dff_q_4)
);
MUX2 mux_inst_2638 (
  .O(mux_o_2638),
  .I0(mux_o_2608),
  .I1(mux_o_2609),
  .S0(dff_q_4)
);
MUX2 mux_inst_2639 (
  .O(mux_o_2639),
  .I0(mux_o_2610),
  .I1(mux_o_2611),
  .S0(dff_q_4)
);
MUX2 mux_inst_2640 (
  .O(mux_o_2640),
  .I0(mux_o_2612),
  .I1(mux_o_2613),
  .S0(dff_q_4)
);
MUX2 mux_inst_2641 (
  .O(mux_o_2641),
  .I0(mux_o_2614),
  .I1(mux_o_2615),
  .S0(dff_q_4)
);
MUX2 mux_inst_2642 (
  .O(mux_o_2642),
  .I0(mux_o_2616),
  .I1(mux_o_2617),
  .S0(dff_q_4)
);
MUX2 mux_inst_2643 (
  .O(mux_o_2643),
  .I0(mux_o_2618),
  .I1(mux_o_2619),
  .S0(dff_q_4)
);
MUX2 mux_inst_2644 (
  .O(mux_o_2644),
  .I0(mux_o_2620),
  .I1(mux_o_2621),
  .S0(dff_q_4)
);
MUX2 mux_inst_2645 (
  .O(mux_o_2645),
  .I0(mux_o_2622),
  .I1(mux_o_2623),
  .S0(dff_q_4)
);
MUX2 mux_inst_2646 (
  .O(mux_o_2646),
  .I0(mux_o_2624),
  .I1(mux_o_2625),
  .S0(dff_q_4)
);
MUX2 mux_inst_2647 (
  .O(mux_o_2647),
  .I0(mux_o_2626),
  .I1(mux_o_2627),
  .S0(dff_q_4)
);
MUX2 mux_inst_2648 (
  .O(mux_o_2648),
  .I0(mux_o_2628),
  .I1(mux_o_2629),
  .S0(dff_q_4)
);
MUX2 mux_inst_2649 (
  .O(mux_o_2649),
  .I0(mux_o_2630),
  .I1(mux_o_2631),
  .S0(dff_q_4)
);
MUX2 mux_inst_2650 (
  .O(mux_o_2650),
  .I0(mux_o_2632),
  .I1(mux_o_2633),
  .S0(dff_q_4)
);
MUX2 mux_inst_2651 (
  .O(mux_o_2651),
  .I0(mux_o_2634),
  .I1(mux_o_2635),
  .S0(dff_q_4)
);
MUX2 mux_inst_2652 (
  .O(mux_o_2652),
  .I0(mux_o_2636),
  .I1(mux_o_2637),
  .S0(dff_q_3)
);
MUX2 mux_inst_2653 (
  .O(mux_o_2653),
  .I0(mux_o_2638),
  .I1(mux_o_2639),
  .S0(dff_q_3)
);
MUX2 mux_inst_2654 (
  .O(mux_o_2654),
  .I0(mux_o_2640),
  .I1(mux_o_2641),
  .S0(dff_q_3)
);
MUX2 mux_inst_2655 (
  .O(mux_o_2655),
  .I0(mux_o_2642),
  .I1(mux_o_2643),
  .S0(dff_q_3)
);
MUX2 mux_inst_2656 (
  .O(mux_o_2656),
  .I0(mux_o_2644),
  .I1(mux_o_2645),
  .S0(dff_q_3)
);
MUX2 mux_inst_2657 (
  .O(mux_o_2657),
  .I0(mux_o_2646),
  .I1(mux_o_2647),
  .S0(dff_q_3)
);
MUX2 mux_inst_2658 (
  .O(mux_o_2658),
  .I0(mux_o_2648),
  .I1(mux_o_2649),
  .S0(dff_q_3)
);
MUX2 mux_inst_2659 (
  .O(mux_o_2659),
  .I0(mux_o_2650),
  .I1(mux_o_2651),
  .S0(dff_q_3)
);
MUX2 mux_inst_2660 (
  .O(mux_o_2660),
  .I0(mux_o_2652),
  .I1(mux_o_2653),
  .S0(dff_q_2)
);
MUX2 mux_inst_2661 (
  .O(mux_o_2661),
  .I0(mux_o_2654),
  .I1(mux_o_2655),
  .S0(dff_q_2)
);
MUX2 mux_inst_2662 (
  .O(mux_o_2662),
  .I0(mux_o_2656),
  .I1(mux_o_2657),
  .S0(dff_q_2)
);
MUX2 mux_inst_2663 (
  .O(mux_o_2663),
  .I0(mux_o_2658),
  .I1(mux_o_2659),
  .S0(dff_q_2)
);
MUX2 mux_inst_2664 (
  .O(mux_o_2664),
  .I0(mux_o_2660),
  .I1(mux_o_2661),
  .S0(dff_q_1)
);
MUX2 mux_inst_2665 (
  .O(mux_o_2665),
  .I0(mux_o_2662),
  .I1(mux_o_2663),
  .S0(dff_q_1)
);
MUX2 mux_inst_2666 (
  .O(dout[20]),
  .I0(mux_o_2664),
  .I1(mux_o_2665),
  .S0(dff_q_0)
);
MUX2 mux_inst_2667 (
  .O(mux_o_2667),
  .I0(sdpb_inst_128_dout[21]),
  .I1(sdpb_inst_129_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2668 (
  .O(mux_o_2668),
  .I0(sdpb_inst_130_dout[21]),
  .I1(sdpb_inst_131_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2669 (
  .O(mux_o_2669),
  .I0(sdpb_inst_132_dout[21]),
  .I1(sdpb_inst_133_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2670 (
  .O(mux_o_2670),
  .I0(sdpb_inst_134_dout[21]),
  .I1(sdpb_inst_135_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2671 (
  .O(mux_o_2671),
  .I0(sdpb_inst_136_dout[21]),
  .I1(sdpb_inst_137_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2672 (
  .O(mux_o_2672),
  .I0(sdpb_inst_138_dout[21]),
  .I1(sdpb_inst_139_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2673 (
  .O(mux_o_2673),
  .I0(sdpb_inst_140_dout[21]),
  .I1(sdpb_inst_141_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2674 (
  .O(mux_o_2674),
  .I0(sdpb_inst_142_dout[21]),
  .I1(sdpb_inst_143_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2675 (
  .O(mux_o_2675),
  .I0(sdpb_inst_144_dout[21]),
  .I1(sdpb_inst_145_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2676 (
  .O(mux_o_2676),
  .I0(sdpb_inst_146_dout[21]),
  .I1(sdpb_inst_147_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2677 (
  .O(mux_o_2677),
  .I0(sdpb_inst_148_dout[21]),
  .I1(sdpb_inst_149_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2678 (
  .O(mux_o_2678),
  .I0(sdpb_inst_150_dout[21]),
  .I1(sdpb_inst_151_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2679 (
  .O(mux_o_2679),
  .I0(sdpb_inst_152_dout[21]),
  .I1(sdpb_inst_153_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2680 (
  .O(mux_o_2680),
  .I0(sdpb_inst_154_dout[21]),
  .I1(sdpb_inst_155_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2681 (
  .O(mux_o_2681),
  .I0(sdpb_inst_156_dout[21]),
  .I1(sdpb_inst_157_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2682 (
  .O(mux_o_2682),
  .I0(sdpb_inst_158_dout[21]),
  .I1(sdpb_inst_159_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2683 (
  .O(mux_o_2683),
  .I0(sdpb_inst_160_dout[21]),
  .I1(sdpb_inst_161_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2684 (
  .O(mux_o_2684),
  .I0(sdpb_inst_162_dout[21]),
  .I1(sdpb_inst_163_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2685 (
  .O(mux_o_2685),
  .I0(sdpb_inst_164_dout[21]),
  .I1(sdpb_inst_165_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2686 (
  .O(mux_o_2686),
  .I0(sdpb_inst_166_dout[21]),
  .I1(sdpb_inst_167_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2687 (
  .O(mux_o_2687),
  .I0(sdpb_inst_168_dout[21]),
  .I1(sdpb_inst_169_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2688 (
  .O(mux_o_2688),
  .I0(sdpb_inst_170_dout[21]),
  .I1(sdpb_inst_171_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2689 (
  .O(mux_o_2689),
  .I0(sdpb_inst_172_dout[21]),
  .I1(sdpb_inst_173_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2690 (
  .O(mux_o_2690),
  .I0(sdpb_inst_174_dout[21]),
  .I1(sdpb_inst_175_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2691 (
  .O(mux_o_2691),
  .I0(sdpb_inst_176_dout[21]),
  .I1(sdpb_inst_177_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2692 (
  .O(mux_o_2692),
  .I0(sdpb_inst_178_dout[21]),
  .I1(sdpb_inst_179_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2693 (
  .O(mux_o_2693),
  .I0(sdpb_inst_180_dout[21]),
  .I1(sdpb_inst_181_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2694 (
  .O(mux_o_2694),
  .I0(sdpb_inst_182_dout[21]),
  .I1(sdpb_inst_183_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2695 (
  .O(mux_o_2695),
  .I0(sdpb_inst_184_dout[21]),
  .I1(sdpb_inst_185_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2696 (
  .O(mux_o_2696),
  .I0(sdpb_inst_186_dout[21]),
  .I1(sdpb_inst_187_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2697 (
  .O(mux_o_2697),
  .I0(sdpb_inst_188_dout[21]),
  .I1(sdpb_inst_189_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2698 (
  .O(mux_o_2698),
  .I0(sdpb_inst_190_dout[21]),
  .I1(sdpb_inst_191_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2699 (
  .O(mux_o_2699),
  .I0(sdpb_inst_192_dout[21]),
  .I1(sdpb_inst_193_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2700 (
  .O(mux_o_2700),
  .I0(sdpb_inst_194_dout[21]),
  .I1(sdpb_inst_195_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2701 (
  .O(mux_o_2701),
  .I0(sdpb_inst_196_dout[21]),
  .I1(sdpb_inst_197_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2702 (
  .O(mux_o_2702),
  .I0(sdpb_inst_198_dout[21]),
  .I1(sdpb_inst_199_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2703 (
  .O(mux_o_2703),
  .I0(sdpb_inst_200_dout[21]),
  .I1(sdpb_inst_201_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2704 (
  .O(mux_o_2704),
  .I0(sdpb_inst_202_dout[21]),
  .I1(sdpb_inst_203_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2705 (
  .O(mux_o_2705),
  .I0(sdpb_inst_204_dout[21]),
  .I1(sdpb_inst_205_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2706 (
  .O(mux_o_2706),
  .I0(sdpb_inst_206_dout[21]),
  .I1(sdpb_inst_207_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2707 (
  .O(mux_o_2707),
  .I0(sdpb_inst_208_dout[21]),
  .I1(sdpb_inst_209_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2708 (
  .O(mux_o_2708),
  .I0(sdpb_inst_210_dout[21]),
  .I1(sdpb_inst_211_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2709 (
  .O(mux_o_2709),
  .I0(sdpb_inst_212_dout[21]),
  .I1(sdpb_inst_213_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2710 (
  .O(mux_o_2710),
  .I0(sdpb_inst_214_dout[21]),
  .I1(sdpb_inst_215_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2711 (
  .O(mux_o_2711),
  .I0(sdpb_inst_216_dout[21]),
  .I1(sdpb_inst_217_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2712 (
  .O(mux_o_2712),
  .I0(sdpb_inst_218_dout[21]),
  .I1(sdpb_inst_219_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2713 (
  .O(mux_o_2713),
  .I0(sdpb_inst_220_dout[21]),
  .I1(sdpb_inst_221_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2714 (
  .O(mux_o_2714),
  .I0(sdpb_inst_222_dout[21]),
  .I1(sdpb_inst_223_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2715 (
  .O(mux_o_2715),
  .I0(sdpb_inst_224_dout[21]),
  .I1(sdpb_inst_225_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2716 (
  .O(mux_o_2716),
  .I0(sdpb_inst_226_dout[21]),
  .I1(sdpb_inst_227_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2717 (
  .O(mux_o_2717),
  .I0(sdpb_inst_228_dout[21]),
  .I1(sdpb_inst_229_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2718 (
  .O(mux_o_2718),
  .I0(sdpb_inst_230_dout[21]),
  .I1(sdpb_inst_231_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2719 (
  .O(mux_o_2719),
  .I0(sdpb_inst_232_dout[21]),
  .I1(sdpb_inst_233_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2720 (
  .O(mux_o_2720),
  .I0(sdpb_inst_234_dout[21]),
  .I1(sdpb_inst_235_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2721 (
  .O(mux_o_2721),
  .I0(sdpb_inst_236_dout[21]),
  .I1(sdpb_inst_237_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2722 (
  .O(mux_o_2722),
  .I0(sdpb_inst_238_dout[21]),
  .I1(sdpb_inst_239_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2723 (
  .O(mux_o_2723),
  .I0(sdpb_inst_240_dout[21]),
  .I1(sdpb_inst_241_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2724 (
  .O(mux_o_2724),
  .I0(sdpb_inst_242_dout[21]),
  .I1(sdpb_inst_243_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2725 (
  .O(mux_o_2725),
  .I0(sdpb_inst_244_dout[21]),
  .I1(sdpb_inst_245_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2726 (
  .O(mux_o_2726),
  .I0(sdpb_inst_246_dout[21]),
  .I1(sdpb_inst_247_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2727 (
  .O(mux_o_2727),
  .I0(sdpb_inst_248_dout[21]),
  .I1(sdpb_inst_249_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2728 (
  .O(mux_o_2728),
  .I0(sdpb_inst_250_dout[21]),
  .I1(sdpb_inst_251_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2729 (
  .O(mux_o_2729),
  .I0(sdpb_inst_252_dout[21]),
  .I1(sdpb_inst_253_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2730 (
  .O(mux_o_2730),
  .I0(sdpb_inst_254_dout[21]),
  .I1(sdpb_inst_255_dout[21]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2731 (
  .O(mux_o_2731),
  .I0(mux_o_2667),
  .I1(mux_o_2668),
  .S0(dff_q_5)
);
MUX2 mux_inst_2732 (
  .O(mux_o_2732),
  .I0(mux_o_2669),
  .I1(mux_o_2670),
  .S0(dff_q_5)
);
MUX2 mux_inst_2733 (
  .O(mux_o_2733),
  .I0(mux_o_2671),
  .I1(mux_o_2672),
  .S0(dff_q_5)
);
MUX2 mux_inst_2734 (
  .O(mux_o_2734),
  .I0(mux_o_2673),
  .I1(mux_o_2674),
  .S0(dff_q_5)
);
MUX2 mux_inst_2735 (
  .O(mux_o_2735),
  .I0(mux_o_2675),
  .I1(mux_o_2676),
  .S0(dff_q_5)
);
MUX2 mux_inst_2736 (
  .O(mux_o_2736),
  .I0(mux_o_2677),
  .I1(mux_o_2678),
  .S0(dff_q_5)
);
MUX2 mux_inst_2737 (
  .O(mux_o_2737),
  .I0(mux_o_2679),
  .I1(mux_o_2680),
  .S0(dff_q_5)
);
MUX2 mux_inst_2738 (
  .O(mux_o_2738),
  .I0(mux_o_2681),
  .I1(mux_o_2682),
  .S0(dff_q_5)
);
MUX2 mux_inst_2739 (
  .O(mux_o_2739),
  .I0(mux_o_2683),
  .I1(mux_o_2684),
  .S0(dff_q_5)
);
MUX2 mux_inst_2740 (
  .O(mux_o_2740),
  .I0(mux_o_2685),
  .I1(mux_o_2686),
  .S0(dff_q_5)
);
MUX2 mux_inst_2741 (
  .O(mux_o_2741),
  .I0(mux_o_2687),
  .I1(mux_o_2688),
  .S0(dff_q_5)
);
MUX2 mux_inst_2742 (
  .O(mux_o_2742),
  .I0(mux_o_2689),
  .I1(mux_o_2690),
  .S0(dff_q_5)
);
MUX2 mux_inst_2743 (
  .O(mux_o_2743),
  .I0(mux_o_2691),
  .I1(mux_o_2692),
  .S0(dff_q_5)
);
MUX2 mux_inst_2744 (
  .O(mux_o_2744),
  .I0(mux_o_2693),
  .I1(mux_o_2694),
  .S0(dff_q_5)
);
MUX2 mux_inst_2745 (
  .O(mux_o_2745),
  .I0(mux_o_2695),
  .I1(mux_o_2696),
  .S0(dff_q_5)
);
MUX2 mux_inst_2746 (
  .O(mux_o_2746),
  .I0(mux_o_2697),
  .I1(mux_o_2698),
  .S0(dff_q_5)
);
MUX2 mux_inst_2747 (
  .O(mux_o_2747),
  .I0(mux_o_2699),
  .I1(mux_o_2700),
  .S0(dff_q_5)
);
MUX2 mux_inst_2748 (
  .O(mux_o_2748),
  .I0(mux_o_2701),
  .I1(mux_o_2702),
  .S0(dff_q_5)
);
MUX2 mux_inst_2749 (
  .O(mux_o_2749),
  .I0(mux_o_2703),
  .I1(mux_o_2704),
  .S0(dff_q_5)
);
MUX2 mux_inst_2750 (
  .O(mux_o_2750),
  .I0(mux_o_2705),
  .I1(mux_o_2706),
  .S0(dff_q_5)
);
MUX2 mux_inst_2751 (
  .O(mux_o_2751),
  .I0(mux_o_2707),
  .I1(mux_o_2708),
  .S0(dff_q_5)
);
MUX2 mux_inst_2752 (
  .O(mux_o_2752),
  .I0(mux_o_2709),
  .I1(mux_o_2710),
  .S0(dff_q_5)
);
MUX2 mux_inst_2753 (
  .O(mux_o_2753),
  .I0(mux_o_2711),
  .I1(mux_o_2712),
  .S0(dff_q_5)
);
MUX2 mux_inst_2754 (
  .O(mux_o_2754),
  .I0(mux_o_2713),
  .I1(mux_o_2714),
  .S0(dff_q_5)
);
MUX2 mux_inst_2755 (
  .O(mux_o_2755),
  .I0(mux_o_2715),
  .I1(mux_o_2716),
  .S0(dff_q_5)
);
MUX2 mux_inst_2756 (
  .O(mux_o_2756),
  .I0(mux_o_2717),
  .I1(mux_o_2718),
  .S0(dff_q_5)
);
MUX2 mux_inst_2757 (
  .O(mux_o_2757),
  .I0(mux_o_2719),
  .I1(mux_o_2720),
  .S0(dff_q_5)
);
MUX2 mux_inst_2758 (
  .O(mux_o_2758),
  .I0(mux_o_2721),
  .I1(mux_o_2722),
  .S0(dff_q_5)
);
MUX2 mux_inst_2759 (
  .O(mux_o_2759),
  .I0(mux_o_2723),
  .I1(mux_o_2724),
  .S0(dff_q_5)
);
MUX2 mux_inst_2760 (
  .O(mux_o_2760),
  .I0(mux_o_2725),
  .I1(mux_o_2726),
  .S0(dff_q_5)
);
MUX2 mux_inst_2761 (
  .O(mux_o_2761),
  .I0(mux_o_2727),
  .I1(mux_o_2728),
  .S0(dff_q_5)
);
MUX2 mux_inst_2762 (
  .O(mux_o_2762),
  .I0(mux_o_2729),
  .I1(mux_o_2730),
  .S0(dff_q_5)
);
MUX2 mux_inst_2763 (
  .O(mux_o_2763),
  .I0(mux_o_2731),
  .I1(mux_o_2732),
  .S0(dff_q_4)
);
MUX2 mux_inst_2764 (
  .O(mux_o_2764),
  .I0(mux_o_2733),
  .I1(mux_o_2734),
  .S0(dff_q_4)
);
MUX2 mux_inst_2765 (
  .O(mux_o_2765),
  .I0(mux_o_2735),
  .I1(mux_o_2736),
  .S0(dff_q_4)
);
MUX2 mux_inst_2766 (
  .O(mux_o_2766),
  .I0(mux_o_2737),
  .I1(mux_o_2738),
  .S0(dff_q_4)
);
MUX2 mux_inst_2767 (
  .O(mux_o_2767),
  .I0(mux_o_2739),
  .I1(mux_o_2740),
  .S0(dff_q_4)
);
MUX2 mux_inst_2768 (
  .O(mux_o_2768),
  .I0(mux_o_2741),
  .I1(mux_o_2742),
  .S0(dff_q_4)
);
MUX2 mux_inst_2769 (
  .O(mux_o_2769),
  .I0(mux_o_2743),
  .I1(mux_o_2744),
  .S0(dff_q_4)
);
MUX2 mux_inst_2770 (
  .O(mux_o_2770),
  .I0(mux_o_2745),
  .I1(mux_o_2746),
  .S0(dff_q_4)
);
MUX2 mux_inst_2771 (
  .O(mux_o_2771),
  .I0(mux_o_2747),
  .I1(mux_o_2748),
  .S0(dff_q_4)
);
MUX2 mux_inst_2772 (
  .O(mux_o_2772),
  .I0(mux_o_2749),
  .I1(mux_o_2750),
  .S0(dff_q_4)
);
MUX2 mux_inst_2773 (
  .O(mux_o_2773),
  .I0(mux_o_2751),
  .I1(mux_o_2752),
  .S0(dff_q_4)
);
MUX2 mux_inst_2774 (
  .O(mux_o_2774),
  .I0(mux_o_2753),
  .I1(mux_o_2754),
  .S0(dff_q_4)
);
MUX2 mux_inst_2775 (
  .O(mux_o_2775),
  .I0(mux_o_2755),
  .I1(mux_o_2756),
  .S0(dff_q_4)
);
MUX2 mux_inst_2776 (
  .O(mux_o_2776),
  .I0(mux_o_2757),
  .I1(mux_o_2758),
  .S0(dff_q_4)
);
MUX2 mux_inst_2777 (
  .O(mux_o_2777),
  .I0(mux_o_2759),
  .I1(mux_o_2760),
  .S0(dff_q_4)
);
MUX2 mux_inst_2778 (
  .O(mux_o_2778),
  .I0(mux_o_2761),
  .I1(mux_o_2762),
  .S0(dff_q_4)
);
MUX2 mux_inst_2779 (
  .O(mux_o_2779),
  .I0(mux_o_2763),
  .I1(mux_o_2764),
  .S0(dff_q_3)
);
MUX2 mux_inst_2780 (
  .O(mux_o_2780),
  .I0(mux_o_2765),
  .I1(mux_o_2766),
  .S0(dff_q_3)
);
MUX2 mux_inst_2781 (
  .O(mux_o_2781),
  .I0(mux_o_2767),
  .I1(mux_o_2768),
  .S0(dff_q_3)
);
MUX2 mux_inst_2782 (
  .O(mux_o_2782),
  .I0(mux_o_2769),
  .I1(mux_o_2770),
  .S0(dff_q_3)
);
MUX2 mux_inst_2783 (
  .O(mux_o_2783),
  .I0(mux_o_2771),
  .I1(mux_o_2772),
  .S0(dff_q_3)
);
MUX2 mux_inst_2784 (
  .O(mux_o_2784),
  .I0(mux_o_2773),
  .I1(mux_o_2774),
  .S0(dff_q_3)
);
MUX2 mux_inst_2785 (
  .O(mux_o_2785),
  .I0(mux_o_2775),
  .I1(mux_o_2776),
  .S0(dff_q_3)
);
MUX2 mux_inst_2786 (
  .O(mux_o_2786),
  .I0(mux_o_2777),
  .I1(mux_o_2778),
  .S0(dff_q_3)
);
MUX2 mux_inst_2787 (
  .O(mux_o_2787),
  .I0(mux_o_2779),
  .I1(mux_o_2780),
  .S0(dff_q_2)
);
MUX2 mux_inst_2788 (
  .O(mux_o_2788),
  .I0(mux_o_2781),
  .I1(mux_o_2782),
  .S0(dff_q_2)
);
MUX2 mux_inst_2789 (
  .O(mux_o_2789),
  .I0(mux_o_2783),
  .I1(mux_o_2784),
  .S0(dff_q_2)
);
MUX2 mux_inst_2790 (
  .O(mux_o_2790),
  .I0(mux_o_2785),
  .I1(mux_o_2786),
  .S0(dff_q_2)
);
MUX2 mux_inst_2791 (
  .O(mux_o_2791),
  .I0(mux_o_2787),
  .I1(mux_o_2788),
  .S0(dff_q_1)
);
MUX2 mux_inst_2792 (
  .O(mux_o_2792),
  .I0(mux_o_2789),
  .I1(mux_o_2790),
  .S0(dff_q_1)
);
MUX2 mux_inst_2793 (
  .O(dout[21]),
  .I0(mux_o_2791),
  .I1(mux_o_2792),
  .S0(dff_q_0)
);
MUX2 mux_inst_2794 (
  .O(mux_o_2794),
  .I0(sdpb_inst_128_dout[22]),
  .I1(sdpb_inst_129_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2795 (
  .O(mux_o_2795),
  .I0(sdpb_inst_130_dout[22]),
  .I1(sdpb_inst_131_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2796 (
  .O(mux_o_2796),
  .I0(sdpb_inst_132_dout[22]),
  .I1(sdpb_inst_133_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2797 (
  .O(mux_o_2797),
  .I0(sdpb_inst_134_dout[22]),
  .I1(sdpb_inst_135_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2798 (
  .O(mux_o_2798),
  .I0(sdpb_inst_136_dout[22]),
  .I1(sdpb_inst_137_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2799 (
  .O(mux_o_2799),
  .I0(sdpb_inst_138_dout[22]),
  .I1(sdpb_inst_139_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2800 (
  .O(mux_o_2800),
  .I0(sdpb_inst_140_dout[22]),
  .I1(sdpb_inst_141_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2801 (
  .O(mux_o_2801),
  .I0(sdpb_inst_142_dout[22]),
  .I1(sdpb_inst_143_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2802 (
  .O(mux_o_2802),
  .I0(sdpb_inst_144_dout[22]),
  .I1(sdpb_inst_145_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2803 (
  .O(mux_o_2803),
  .I0(sdpb_inst_146_dout[22]),
  .I1(sdpb_inst_147_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2804 (
  .O(mux_o_2804),
  .I0(sdpb_inst_148_dout[22]),
  .I1(sdpb_inst_149_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2805 (
  .O(mux_o_2805),
  .I0(sdpb_inst_150_dout[22]),
  .I1(sdpb_inst_151_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2806 (
  .O(mux_o_2806),
  .I0(sdpb_inst_152_dout[22]),
  .I1(sdpb_inst_153_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2807 (
  .O(mux_o_2807),
  .I0(sdpb_inst_154_dout[22]),
  .I1(sdpb_inst_155_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2808 (
  .O(mux_o_2808),
  .I0(sdpb_inst_156_dout[22]),
  .I1(sdpb_inst_157_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2809 (
  .O(mux_o_2809),
  .I0(sdpb_inst_158_dout[22]),
  .I1(sdpb_inst_159_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2810 (
  .O(mux_o_2810),
  .I0(sdpb_inst_160_dout[22]),
  .I1(sdpb_inst_161_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2811 (
  .O(mux_o_2811),
  .I0(sdpb_inst_162_dout[22]),
  .I1(sdpb_inst_163_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2812 (
  .O(mux_o_2812),
  .I0(sdpb_inst_164_dout[22]),
  .I1(sdpb_inst_165_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2813 (
  .O(mux_o_2813),
  .I0(sdpb_inst_166_dout[22]),
  .I1(sdpb_inst_167_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2814 (
  .O(mux_o_2814),
  .I0(sdpb_inst_168_dout[22]),
  .I1(sdpb_inst_169_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2815 (
  .O(mux_o_2815),
  .I0(sdpb_inst_170_dout[22]),
  .I1(sdpb_inst_171_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2816 (
  .O(mux_o_2816),
  .I0(sdpb_inst_172_dout[22]),
  .I1(sdpb_inst_173_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2817 (
  .O(mux_o_2817),
  .I0(sdpb_inst_174_dout[22]),
  .I1(sdpb_inst_175_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2818 (
  .O(mux_o_2818),
  .I0(sdpb_inst_176_dout[22]),
  .I1(sdpb_inst_177_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2819 (
  .O(mux_o_2819),
  .I0(sdpb_inst_178_dout[22]),
  .I1(sdpb_inst_179_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2820 (
  .O(mux_o_2820),
  .I0(sdpb_inst_180_dout[22]),
  .I1(sdpb_inst_181_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2821 (
  .O(mux_o_2821),
  .I0(sdpb_inst_182_dout[22]),
  .I1(sdpb_inst_183_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2822 (
  .O(mux_o_2822),
  .I0(sdpb_inst_184_dout[22]),
  .I1(sdpb_inst_185_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2823 (
  .O(mux_o_2823),
  .I0(sdpb_inst_186_dout[22]),
  .I1(sdpb_inst_187_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2824 (
  .O(mux_o_2824),
  .I0(sdpb_inst_188_dout[22]),
  .I1(sdpb_inst_189_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2825 (
  .O(mux_o_2825),
  .I0(sdpb_inst_190_dout[22]),
  .I1(sdpb_inst_191_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2826 (
  .O(mux_o_2826),
  .I0(sdpb_inst_192_dout[22]),
  .I1(sdpb_inst_193_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2827 (
  .O(mux_o_2827),
  .I0(sdpb_inst_194_dout[22]),
  .I1(sdpb_inst_195_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2828 (
  .O(mux_o_2828),
  .I0(sdpb_inst_196_dout[22]),
  .I1(sdpb_inst_197_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2829 (
  .O(mux_o_2829),
  .I0(sdpb_inst_198_dout[22]),
  .I1(sdpb_inst_199_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2830 (
  .O(mux_o_2830),
  .I0(sdpb_inst_200_dout[22]),
  .I1(sdpb_inst_201_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2831 (
  .O(mux_o_2831),
  .I0(sdpb_inst_202_dout[22]),
  .I1(sdpb_inst_203_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2832 (
  .O(mux_o_2832),
  .I0(sdpb_inst_204_dout[22]),
  .I1(sdpb_inst_205_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2833 (
  .O(mux_o_2833),
  .I0(sdpb_inst_206_dout[22]),
  .I1(sdpb_inst_207_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2834 (
  .O(mux_o_2834),
  .I0(sdpb_inst_208_dout[22]),
  .I1(sdpb_inst_209_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2835 (
  .O(mux_o_2835),
  .I0(sdpb_inst_210_dout[22]),
  .I1(sdpb_inst_211_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2836 (
  .O(mux_o_2836),
  .I0(sdpb_inst_212_dout[22]),
  .I1(sdpb_inst_213_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2837 (
  .O(mux_o_2837),
  .I0(sdpb_inst_214_dout[22]),
  .I1(sdpb_inst_215_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2838 (
  .O(mux_o_2838),
  .I0(sdpb_inst_216_dout[22]),
  .I1(sdpb_inst_217_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2839 (
  .O(mux_o_2839),
  .I0(sdpb_inst_218_dout[22]),
  .I1(sdpb_inst_219_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2840 (
  .O(mux_o_2840),
  .I0(sdpb_inst_220_dout[22]),
  .I1(sdpb_inst_221_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2841 (
  .O(mux_o_2841),
  .I0(sdpb_inst_222_dout[22]),
  .I1(sdpb_inst_223_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2842 (
  .O(mux_o_2842),
  .I0(sdpb_inst_224_dout[22]),
  .I1(sdpb_inst_225_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2843 (
  .O(mux_o_2843),
  .I0(sdpb_inst_226_dout[22]),
  .I1(sdpb_inst_227_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2844 (
  .O(mux_o_2844),
  .I0(sdpb_inst_228_dout[22]),
  .I1(sdpb_inst_229_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2845 (
  .O(mux_o_2845),
  .I0(sdpb_inst_230_dout[22]),
  .I1(sdpb_inst_231_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2846 (
  .O(mux_o_2846),
  .I0(sdpb_inst_232_dout[22]),
  .I1(sdpb_inst_233_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2847 (
  .O(mux_o_2847),
  .I0(sdpb_inst_234_dout[22]),
  .I1(sdpb_inst_235_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2848 (
  .O(mux_o_2848),
  .I0(sdpb_inst_236_dout[22]),
  .I1(sdpb_inst_237_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2849 (
  .O(mux_o_2849),
  .I0(sdpb_inst_238_dout[22]),
  .I1(sdpb_inst_239_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2850 (
  .O(mux_o_2850),
  .I0(sdpb_inst_240_dout[22]),
  .I1(sdpb_inst_241_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2851 (
  .O(mux_o_2851),
  .I0(sdpb_inst_242_dout[22]),
  .I1(sdpb_inst_243_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2852 (
  .O(mux_o_2852),
  .I0(sdpb_inst_244_dout[22]),
  .I1(sdpb_inst_245_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2853 (
  .O(mux_o_2853),
  .I0(sdpb_inst_246_dout[22]),
  .I1(sdpb_inst_247_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2854 (
  .O(mux_o_2854),
  .I0(sdpb_inst_248_dout[22]),
  .I1(sdpb_inst_249_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2855 (
  .O(mux_o_2855),
  .I0(sdpb_inst_250_dout[22]),
  .I1(sdpb_inst_251_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2856 (
  .O(mux_o_2856),
  .I0(sdpb_inst_252_dout[22]),
  .I1(sdpb_inst_253_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2857 (
  .O(mux_o_2857),
  .I0(sdpb_inst_254_dout[22]),
  .I1(sdpb_inst_255_dout[22]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2858 (
  .O(mux_o_2858),
  .I0(mux_o_2794),
  .I1(mux_o_2795),
  .S0(dff_q_5)
);
MUX2 mux_inst_2859 (
  .O(mux_o_2859),
  .I0(mux_o_2796),
  .I1(mux_o_2797),
  .S0(dff_q_5)
);
MUX2 mux_inst_2860 (
  .O(mux_o_2860),
  .I0(mux_o_2798),
  .I1(mux_o_2799),
  .S0(dff_q_5)
);
MUX2 mux_inst_2861 (
  .O(mux_o_2861),
  .I0(mux_o_2800),
  .I1(mux_o_2801),
  .S0(dff_q_5)
);
MUX2 mux_inst_2862 (
  .O(mux_o_2862),
  .I0(mux_o_2802),
  .I1(mux_o_2803),
  .S0(dff_q_5)
);
MUX2 mux_inst_2863 (
  .O(mux_o_2863),
  .I0(mux_o_2804),
  .I1(mux_o_2805),
  .S0(dff_q_5)
);
MUX2 mux_inst_2864 (
  .O(mux_o_2864),
  .I0(mux_o_2806),
  .I1(mux_o_2807),
  .S0(dff_q_5)
);
MUX2 mux_inst_2865 (
  .O(mux_o_2865),
  .I0(mux_o_2808),
  .I1(mux_o_2809),
  .S0(dff_q_5)
);
MUX2 mux_inst_2866 (
  .O(mux_o_2866),
  .I0(mux_o_2810),
  .I1(mux_o_2811),
  .S0(dff_q_5)
);
MUX2 mux_inst_2867 (
  .O(mux_o_2867),
  .I0(mux_o_2812),
  .I1(mux_o_2813),
  .S0(dff_q_5)
);
MUX2 mux_inst_2868 (
  .O(mux_o_2868),
  .I0(mux_o_2814),
  .I1(mux_o_2815),
  .S0(dff_q_5)
);
MUX2 mux_inst_2869 (
  .O(mux_o_2869),
  .I0(mux_o_2816),
  .I1(mux_o_2817),
  .S0(dff_q_5)
);
MUX2 mux_inst_2870 (
  .O(mux_o_2870),
  .I0(mux_o_2818),
  .I1(mux_o_2819),
  .S0(dff_q_5)
);
MUX2 mux_inst_2871 (
  .O(mux_o_2871),
  .I0(mux_o_2820),
  .I1(mux_o_2821),
  .S0(dff_q_5)
);
MUX2 mux_inst_2872 (
  .O(mux_o_2872),
  .I0(mux_o_2822),
  .I1(mux_o_2823),
  .S0(dff_q_5)
);
MUX2 mux_inst_2873 (
  .O(mux_o_2873),
  .I0(mux_o_2824),
  .I1(mux_o_2825),
  .S0(dff_q_5)
);
MUX2 mux_inst_2874 (
  .O(mux_o_2874),
  .I0(mux_o_2826),
  .I1(mux_o_2827),
  .S0(dff_q_5)
);
MUX2 mux_inst_2875 (
  .O(mux_o_2875),
  .I0(mux_o_2828),
  .I1(mux_o_2829),
  .S0(dff_q_5)
);
MUX2 mux_inst_2876 (
  .O(mux_o_2876),
  .I0(mux_o_2830),
  .I1(mux_o_2831),
  .S0(dff_q_5)
);
MUX2 mux_inst_2877 (
  .O(mux_o_2877),
  .I0(mux_o_2832),
  .I1(mux_o_2833),
  .S0(dff_q_5)
);
MUX2 mux_inst_2878 (
  .O(mux_o_2878),
  .I0(mux_o_2834),
  .I1(mux_o_2835),
  .S0(dff_q_5)
);
MUX2 mux_inst_2879 (
  .O(mux_o_2879),
  .I0(mux_o_2836),
  .I1(mux_o_2837),
  .S0(dff_q_5)
);
MUX2 mux_inst_2880 (
  .O(mux_o_2880),
  .I0(mux_o_2838),
  .I1(mux_o_2839),
  .S0(dff_q_5)
);
MUX2 mux_inst_2881 (
  .O(mux_o_2881),
  .I0(mux_o_2840),
  .I1(mux_o_2841),
  .S0(dff_q_5)
);
MUX2 mux_inst_2882 (
  .O(mux_o_2882),
  .I0(mux_o_2842),
  .I1(mux_o_2843),
  .S0(dff_q_5)
);
MUX2 mux_inst_2883 (
  .O(mux_o_2883),
  .I0(mux_o_2844),
  .I1(mux_o_2845),
  .S0(dff_q_5)
);
MUX2 mux_inst_2884 (
  .O(mux_o_2884),
  .I0(mux_o_2846),
  .I1(mux_o_2847),
  .S0(dff_q_5)
);
MUX2 mux_inst_2885 (
  .O(mux_o_2885),
  .I0(mux_o_2848),
  .I1(mux_o_2849),
  .S0(dff_q_5)
);
MUX2 mux_inst_2886 (
  .O(mux_o_2886),
  .I0(mux_o_2850),
  .I1(mux_o_2851),
  .S0(dff_q_5)
);
MUX2 mux_inst_2887 (
  .O(mux_o_2887),
  .I0(mux_o_2852),
  .I1(mux_o_2853),
  .S0(dff_q_5)
);
MUX2 mux_inst_2888 (
  .O(mux_o_2888),
  .I0(mux_o_2854),
  .I1(mux_o_2855),
  .S0(dff_q_5)
);
MUX2 mux_inst_2889 (
  .O(mux_o_2889),
  .I0(mux_o_2856),
  .I1(mux_o_2857),
  .S0(dff_q_5)
);
MUX2 mux_inst_2890 (
  .O(mux_o_2890),
  .I0(mux_o_2858),
  .I1(mux_o_2859),
  .S0(dff_q_4)
);
MUX2 mux_inst_2891 (
  .O(mux_o_2891),
  .I0(mux_o_2860),
  .I1(mux_o_2861),
  .S0(dff_q_4)
);
MUX2 mux_inst_2892 (
  .O(mux_o_2892),
  .I0(mux_o_2862),
  .I1(mux_o_2863),
  .S0(dff_q_4)
);
MUX2 mux_inst_2893 (
  .O(mux_o_2893),
  .I0(mux_o_2864),
  .I1(mux_o_2865),
  .S0(dff_q_4)
);
MUX2 mux_inst_2894 (
  .O(mux_o_2894),
  .I0(mux_o_2866),
  .I1(mux_o_2867),
  .S0(dff_q_4)
);
MUX2 mux_inst_2895 (
  .O(mux_o_2895),
  .I0(mux_o_2868),
  .I1(mux_o_2869),
  .S0(dff_q_4)
);
MUX2 mux_inst_2896 (
  .O(mux_o_2896),
  .I0(mux_o_2870),
  .I1(mux_o_2871),
  .S0(dff_q_4)
);
MUX2 mux_inst_2897 (
  .O(mux_o_2897),
  .I0(mux_o_2872),
  .I1(mux_o_2873),
  .S0(dff_q_4)
);
MUX2 mux_inst_2898 (
  .O(mux_o_2898),
  .I0(mux_o_2874),
  .I1(mux_o_2875),
  .S0(dff_q_4)
);
MUX2 mux_inst_2899 (
  .O(mux_o_2899),
  .I0(mux_o_2876),
  .I1(mux_o_2877),
  .S0(dff_q_4)
);
MUX2 mux_inst_2900 (
  .O(mux_o_2900),
  .I0(mux_o_2878),
  .I1(mux_o_2879),
  .S0(dff_q_4)
);
MUX2 mux_inst_2901 (
  .O(mux_o_2901),
  .I0(mux_o_2880),
  .I1(mux_o_2881),
  .S0(dff_q_4)
);
MUX2 mux_inst_2902 (
  .O(mux_o_2902),
  .I0(mux_o_2882),
  .I1(mux_o_2883),
  .S0(dff_q_4)
);
MUX2 mux_inst_2903 (
  .O(mux_o_2903),
  .I0(mux_o_2884),
  .I1(mux_o_2885),
  .S0(dff_q_4)
);
MUX2 mux_inst_2904 (
  .O(mux_o_2904),
  .I0(mux_o_2886),
  .I1(mux_o_2887),
  .S0(dff_q_4)
);
MUX2 mux_inst_2905 (
  .O(mux_o_2905),
  .I0(mux_o_2888),
  .I1(mux_o_2889),
  .S0(dff_q_4)
);
MUX2 mux_inst_2906 (
  .O(mux_o_2906),
  .I0(mux_o_2890),
  .I1(mux_o_2891),
  .S0(dff_q_3)
);
MUX2 mux_inst_2907 (
  .O(mux_o_2907),
  .I0(mux_o_2892),
  .I1(mux_o_2893),
  .S0(dff_q_3)
);
MUX2 mux_inst_2908 (
  .O(mux_o_2908),
  .I0(mux_o_2894),
  .I1(mux_o_2895),
  .S0(dff_q_3)
);
MUX2 mux_inst_2909 (
  .O(mux_o_2909),
  .I0(mux_o_2896),
  .I1(mux_o_2897),
  .S0(dff_q_3)
);
MUX2 mux_inst_2910 (
  .O(mux_o_2910),
  .I0(mux_o_2898),
  .I1(mux_o_2899),
  .S0(dff_q_3)
);
MUX2 mux_inst_2911 (
  .O(mux_o_2911),
  .I0(mux_o_2900),
  .I1(mux_o_2901),
  .S0(dff_q_3)
);
MUX2 mux_inst_2912 (
  .O(mux_o_2912),
  .I0(mux_o_2902),
  .I1(mux_o_2903),
  .S0(dff_q_3)
);
MUX2 mux_inst_2913 (
  .O(mux_o_2913),
  .I0(mux_o_2904),
  .I1(mux_o_2905),
  .S0(dff_q_3)
);
MUX2 mux_inst_2914 (
  .O(mux_o_2914),
  .I0(mux_o_2906),
  .I1(mux_o_2907),
  .S0(dff_q_2)
);
MUX2 mux_inst_2915 (
  .O(mux_o_2915),
  .I0(mux_o_2908),
  .I1(mux_o_2909),
  .S0(dff_q_2)
);
MUX2 mux_inst_2916 (
  .O(mux_o_2916),
  .I0(mux_o_2910),
  .I1(mux_o_2911),
  .S0(dff_q_2)
);
MUX2 mux_inst_2917 (
  .O(mux_o_2917),
  .I0(mux_o_2912),
  .I1(mux_o_2913),
  .S0(dff_q_2)
);
MUX2 mux_inst_2918 (
  .O(mux_o_2918),
  .I0(mux_o_2914),
  .I1(mux_o_2915),
  .S0(dff_q_1)
);
MUX2 mux_inst_2919 (
  .O(mux_o_2919),
  .I0(mux_o_2916),
  .I1(mux_o_2917),
  .S0(dff_q_1)
);
MUX2 mux_inst_2920 (
  .O(dout[22]),
  .I0(mux_o_2918),
  .I1(mux_o_2919),
  .S0(dff_q_0)
);
MUX2 mux_inst_2921 (
  .O(mux_o_2921),
  .I0(sdpb_inst_128_dout[23]),
  .I1(sdpb_inst_129_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2922 (
  .O(mux_o_2922),
  .I0(sdpb_inst_130_dout[23]),
  .I1(sdpb_inst_131_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2923 (
  .O(mux_o_2923),
  .I0(sdpb_inst_132_dout[23]),
  .I1(sdpb_inst_133_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2924 (
  .O(mux_o_2924),
  .I0(sdpb_inst_134_dout[23]),
  .I1(sdpb_inst_135_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2925 (
  .O(mux_o_2925),
  .I0(sdpb_inst_136_dout[23]),
  .I1(sdpb_inst_137_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2926 (
  .O(mux_o_2926),
  .I0(sdpb_inst_138_dout[23]),
  .I1(sdpb_inst_139_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2927 (
  .O(mux_o_2927),
  .I0(sdpb_inst_140_dout[23]),
  .I1(sdpb_inst_141_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2928 (
  .O(mux_o_2928),
  .I0(sdpb_inst_142_dout[23]),
  .I1(sdpb_inst_143_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2929 (
  .O(mux_o_2929),
  .I0(sdpb_inst_144_dout[23]),
  .I1(sdpb_inst_145_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2930 (
  .O(mux_o_2930),
  .I0(sdpb_inst_146_dout[23]),
  .I1(sdpb_inst_147_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2931 (
  .O(mux_o_2931),
  .I0(sdpb_inst_148_dout[23]),
  .I1(sdpb_inst_149_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2932 (
  .O(mux_o_2932),
  .I0(sdpb_inst_150_dout[23]),
  .I1(sdpb_inst_151_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2933 (
  .O(mux_o_2933),
  .I0(sdpb_inst_152_dout[23]),
  .I1(sdpb_inst_153_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2934 (
  .O(mux_o_2934),
  .I0(sdpb_inst_154_dout[23]),
  .I1(sdpb_inst_155_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2935 (
  .O(mux_o_2935),
  .I0(sdpb_inst_156_dout[23]),
  .I1(sdpb_inst_157_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2936 (
  .O(mux_o_2936),
  .I0(sdpb_inst_158_dout[23]),
  .I1(sdpb_inst_159_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2937 (
  .O(mux_o_2937),
  .I0(sdpb_inst_160_dout[23]),
  .I1(sdpb_inst_161_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2938 (
  .O(mux_o_2938),
  .I0(sdpb_inst_162_dout[23]),
  .I1(sdpb_inst_163_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2939 (
  .O(mux_o_2939),
  .I0(sdpb_inst_164_dout[23]),
  .I1(sdpb_inst_165_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2940 (
  .O(mux_o_2940),
  .I0(sdpb_inst_166_dout[23]),
  .I1(sdpb_inst_167_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2941 (
  .O(mux_o_2941),
  .I0(sdpb_inst_168_dout[23]),
  .I1(sdpb_inst_169_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2942 (
  .O(mux_o_2942),
  .I0(sdpb_inst_170_dout[23]),
  .I1(sdpb_inst_171_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2943 (
  .O(mux_o_2943),
  .I0(sdpb_inst_172_dout[23]),
  .I1(sdpb_inst_173_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2944 (
  .O(mux_o_2944),
  .I0(sdpb_inst_174_dout[23]),
  .I1(sdpb_inst_175_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2945 (
  .O(mux_o_2945),
  .I0(sdpb_inst_176_dout[23]),
  .I1(sdpb_inst_177_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2946 (
  .O(mux_o_2946),
  .I0(sdpb_inst_178_dout[23]),
  .I1(sdpb_inst_179_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2947 (
  .O(mux_o_2947),
  .I0(sdpb_inst_180_dout[23]),
  .I1(sdpb_inst_181_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2948 (
  .O(mux_o_2948),
  .I0(sdpb_inst_182_dout[23]),
  .I1(sdpb_inst_183_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2949 (
  .O(mux_o_2949),
  .I0(sdpb_inst_184_dout[23]),
  .I1(sdpb_inst_185_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2950 (
  .O(mux_o_2950),
  .I0(sdpb_inst_186_dout[23]),
  .I1(sdpb_inst_187_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2951 (
  .O(mux_o_2951),
  .I0(sdpb_inst_188_dout[23]),
  .I1(sdpb_inst_189_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2952 (
  .O(mux_o_2952),
  .I0(sdpb_inst_190_dout[23]),
  .I1(sdpb_inst_191_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2953 (
  .O(mux_o_2953),
  .I0(sdpb_inst_192_dout[23]),
  .I1(sdpb_inst_193_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2954 (
  .O(mux_o_2954),
  .I0(sdpb_inst_194_dout[23]),
  .I1(sdpb_inst_195_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2955 (
  .O(mux_o_2955),
  .I0(sdpb_inst_196_dout[23]),
  .I1(sdpb_inst_197_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2956 (
  .O(mux_o_2956),
  .I0(sdpb_inst_198_dout[23]),
  .I1(sdpb_inst_199_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2957 (
  .O(mux_o_2957),
  .I0(sdpb_inst_200_dout[23]),
  .I1(sdpb_inst_201_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2958 (
  .O(mux_o_2958),
  .I0(sdpb_inst_202_dout[23]),
  .I1(sdpb_inst_203_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2959 (
  .O(mux_o_2959),
  .I0(sdpb_inst_204_dout[23]),
  .I1(sdpb_inst_205_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2960 (
  .O(mux_o_2960),
  .I0(sdpb_inst_206_dout[23]),
  .I1(sdpb_inst_207_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2961 (
  .O(mux_o_2961),
  .I0(sdpb_inst_208_dout[23]),
  .I1(sdpb_inst_209_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2962 (
  .O(mux_o_2962),
  .I0(sdpb_inst_210_dout[23]),
  .I1(sdpb_inst_211_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2963 (
  .O(mux_o_2963),
  .I0(sdpb_inst_212_dout[23]),
  .I1(sdpb_inst_213_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2964 (
  .O(mux_o_2964),
  .I0(sdpb_inst_214_dout[23]),
  .I1(sdpb_inst_215_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2965 (
  .O(mux_o_2965),
  .I0(sdpb_inst_216_dout[23]),
  .I1(sdpb_inst_217_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2966 (
  .O(mux_o_2966),
  .I0(sdpb_inst_218_dout[23]),
  .I1(sdpb_inst_219_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2967 (
  .O(mux_o_2967),
  .I0(sdpb_inst_220_dout[23]),
  .I1(sdpb_inst_221_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2968 (
  .O(mux_o_2968),
  .I0(sdpb_inst_222_dout[23]),
  .I1(sdpb_inst_223_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2969 (
  .O(mux_o_2969),
  .I0(sdpb_inst_224_dout[23]),
  .I1(sdpb_inst_225_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2970 (
  .O(mux_o_2970),
  .I0(sdpb_inst_226_dout[23]),
  .I1(sdpb_inst_227_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2971 (
  .O(mux_o_2971),
  .I0(sdpb_inst_228_dout[23]),
  .I1(sdpb_inst_229_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2972 (
  .O(mux_o_2972),
  .I0(sdpb_inst_230_dout[23]),
  .I1(sdpb_inst_231_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2973 (
  .O(mux_o_2973),
  .I0(sdpb_inst_232_dout[23]),
  .I1(sdpb_inst_233_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2974 (
  .O(mux_o_2974),
  .I0(sdpb_inst_234_dout[23]),
  .I1(sdpb_inst_235_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2975 (
  .O(mux_o_2975),
  .I0(sdpb_inst_236_dout[23]),
  .I1(sdpb_inst_237_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2976 (
  .O(mux_o_2976),
  .I0(sdpb_inst_238_dout[23]),
  .I1(sdpb_inst_239_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2977 (
  .O(mux_o_2977),
  .I0(sdpb_inst_240_dout[23]),
  .I1(sdpb_inst_241_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2978 (
  .O(mux_o_2978),
  .I0(sdpb_inst_242_dout[23]),
  .I1(sdpb_inst_243_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2979 (
  .O(mux_o_2979),
  .I0(sdpb_inst_244_dout[23]),
  .I1(sdpb_inst_245_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2980 (
  .O(mux_o_2980),
  .I0(sdpb_inst_246_dout[23]),
  .I1(sdpb_inst_247_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2981 (
  .O(mux_o_2981),
  .I0(sdpb_inst_248_dout[23]),
  .I1(sdpb_inst_249_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2982 (
  .O(mux_o_2982),
  .I0(sdpb_inst_250_dout[23]),
  .I1(sdpb_inst_251_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2983 (
  .O(mux_o_2983),
  .I0(sdpb_inst_252_dout[23]),
  .I1(sdpb_inst_253_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2984 (
  .O(mux_o_2984),
  .I0(sdpb_inst_254_dout[23]),
  .I1(sdpb_inst_255_dout[23]),
  .S0(dff_q_6)
);
MUX2 mux_inst_2985 (
  .O(mux_o_2985),
  .I0(mux_o_2921),
  .I1(mux_o_2922),
  .S0(dff_q_5)
);
MUX2 mux_inst_2986 (
  .O(mux_o_2986),
  .I0(mux_o_2923),
  .I1(mux_o_2924),
  .S0(dff_q_5)
);
MUX2 mux_inst_2987 (
  .O(mux_o_2987),
  .I0(mux_o_2925),
  .I1(mux_o_2926),
  .S0(dff_q_5)
);
MUX2 mux_inst_2988 (
  .O(mux_o_2988),
  .I0(mux_o_2927),
  .I1(mux_o_2928),
  .S0(dff_q_5)
);
MUX2 mux_inst_2989 (
  .O(mux_o_2989),
  .I0(mux_o_2929),
  .I1(mux_o_2930),
  .S0(dff_q_5)
);
MUX2 mux_inst_2990 (
  .O(mux_o_2990),
  .I0(mux_o_2931),
  .I1(mux_o_2932),
  .S0(dff_q_5)
);
MUX2 mux_inst_2991 (
  .O(mux_o_2991),
  .I0(mux_o_2933),
  .I1(mux_o_2934),
  .S0(dff_q_5)
);
MUX2 mux_inst_2992 (
  .O(mux_o_2992),
  .I0(mux_o_2935),
  .I1(mux_o_2936),
  .S0(dff_q_5)
);
MUX2 mux_inst_2993 (
  .O(mux_o_2993),
  .I0(mux_o_2937),
  .I1(mux_o_2938),
  .S0(dff_q_5)
);
MUX2 mux_inst_2994 (
  .O(mux_o_2994),
  .I0(mux_o_2939),
  .I1(mux_o_2940),
  .S0(dff_q_5)
);
MUX2 mux_inst_2995 (
  .O(mux_o_2995),
  .I0(mux_o_2941),
  .I1(mux_o_2942),
  .S0(dff_q_5)
);
MUX2 mux_inst_2996 (
  .O(mux_o_2996),
  .I0(mux_o_2943),
  .I1(mux_o_2944),
  .S0(dff_q_5)
);
MUX2 mux_inst_2997 (
  .O(mux_o_2997),
  .I0(mux_o_2945),
  .I1(mux_o_2946),
  .S0(dff_q_5)
);
MUX2 mux_inst_2998 (
  .O(mux_o_2998),
  .I0(mux_o_2947),
  .I1(mux_o_2948),
  .S0(dff_q_5)
);
MUX2 mux_inst_2999 (
  .O(mux_o_2999),
  .I0(mux_o_2949),
  .I1(mux_o_2950),
  .S0(dff_q_5)
);
MUX2 mux_inst_3000 (
  .O(mux_o_3000),
  .I0(mux_o_2951),
  .I1(mux_o_2952),
  .S0(dff_q_5)
);
MUX2 mux_inst_3001 (
  .O(mux_o_3001),
  .I0(mux_o_2953),
  .I1(mux_o_2954),
  .S0(dff_q_5)
);
MUX2 mux_inst_3002 (
  .O(mux_o_3002),
  .I0(mux_o_2955),
  .I1(mux_o_2956),
  .S0(dff_q_5)
);
MUX2 mux_inst_3003 (
  .O(mux_o_3003),
  .I0(mux_o_2957),
  .I1(mux_o_2958),
  .S0(dff_q_5)
);
MUX2 mux_inst_3004 (
  .O(mux_o_3004),
  .I0(mux_o_2959),
  .I1(mux_o_2960),
  .S0(dff_q_5)
);
MUX2 mux_inst_3005 (
  .O(mux_o_3005),
  .I0(mux_o_2961),
  .I1(mux_o_2962),
  .S0(dff_q_5)
);
MUX2 mux_inst_3006 (
  .O(mux_o_3006),
  .I0(mux_o_2963),
  .I1(mux_o_2964),
  .S0(dff_q_5)
);
MUX2 mux_inst_3007 (
  .O(mux_o_3007),
  .I0(mux_o_2965),
  .I1(mux_o_2966),
  .S0(dff_q_5)
);
MUX2 mux_inst_3008 (
  .O(mux_o_3008),
  .I0(mux_o_2967),
  .I1(mux_o_2968),
  .S0(dff_q_5)
);
MUX2 mux_inst_3009 (
  .O(mux_o_3009),
  .I0(mux_o_2969),
  .I1(mux_o_2970),
  .S0(dff_q_5)
);
MUX2 mux_inst_3010 (
  .O(mux_o_3010),
  .I0(mux_o_2971),
  .I1(mux_o_2972),
  .S0(dff_q_5)
);
MUX2 mux_inst_3011 (
  .O(mux_o_3011),
  .I0(mux_o_2973),
  .I1(mux_o_2974),
  .S0(dff_q_5)
);
MUX2 mux_inst_3012 (
  .O(mux_o_3012),
  .I0(mux_o_2975),
  .I1(mux_o_2976),
  .S0(dff_q_5)
);
MUX2 mux_inst_3013 (
  .O(mux_o_3013),
  .I0(mux_o_2977),
  .I1(mux_o_2978),
  .S0(dff_q_5)
);
MUX2 mux_inst_3014 (
  .O(mux_o_3014),
  .I0(mux_o_2979),
  .I1(mux_o_2980),
  .S0(dff_q_5)
);
MUX2 mux_inst_3015 (
  .O(mux_o_3015),
  .I0(mux_o_2981),
  .I1(mux_o_2982),
  .S0(dff_q_5)
);
MUX2 mux_inst_3016 (
  .O(mux_o_3016),
  .I0(mux_o_2983),
  .I1(mux_o_2984),
  .S0(dff_q_5)
);
MUX2 mux_inst_3017 (
  .O(mux_o_3017),
  .I0(mux_o_2985),
  .I1(mux_o_2986),
  .S0(dff_q_4)
);
MUX2 mux_inst_3018 (
  .O(mux_o_3018),
  .I0(mux_o_2987),
  .I1(mux_o_2988),
  .S0(dff_q_4)
);
MUX2 mux_inst_3019 (
  .O(mux_o_3019),
  .I0(mux_o_2989),
  .I1(mux_o_2990),
  .S0(dff_q_4)
);
MUX2 mux_inst_3020 (
  .O(mux_o_3020),
  .I0(mux_o_2991),
  .I1(mux_o_2992),
  .S0(dff_q_4)
);
MUX2 mux_inst_3021 (
  .O(mux_o_3021),
  .I0(mux_o_2993),
  .I1(mux_o_2994),
  .S0(dff_q_4)
);
MUX2 mux_inst_3022 (
  .O(mux_o_3022),
  .I0(mux_o_2995),
  .I1(mux_o_2996),
  .S0(dff_q_4)
);
MUX2 mux_inst_3023 (
  .O(mux_o_3023),
  .I0(mux_o_2997),
  .I1(mux_o_2998),
  .S0(dff_q_4)
);
MUX2 mux_inst_3024 (
  .O(mux_o_3024),
  .I0(mux_o_2999),
  .I1(mux_o_3000),
  .S0(dff_q_4)
);
MUX2 mux_inst_3025 (
  .O(mux_o_3025),
  .I0(mux_o_3001),
  .I1(mux_o_3002),
  .S0(dff_q_4)
);
MUX2 mux_inst_3026 (
  .O(mux_o_3026),
  .I0(mux_o_3003),
  .I1(mux_o_3004),
  .S0(dff_q_4)
);
MUX2 mux_inst_3027 (
  .O(mux_o_3027),
  .I0(mux_o_3005),
  .I1(mux_o_3006),
  .S0(dff_q_4)
);
MUX2 mux_inst_3028 (
  .O(mux_o_3028),
  .I0(mux_o_3007),
  .I1(mux_o_3008),
  .S0(dff_q_4)
);
MUX2 mux_inst_3029 (
  .O(mux_o_3029),
  .I0(mux_o_3009),
  .I1(mux_o_3010),
  .S0(dff_q_4)
);
MUX2 mux_inst_3030 (
  .O(mux_o_3030),
  .I0(mux_o_3011),
  .I1(mux_o_3012),
  .S0(dff_q_4)
);
MUX2 mux_inst_3031 (
  .O(mux_o_3031),
  .I0(mux_o_3013),
  .I1(mux_o_3014),
  .S0(dff_q_4)
);
MUX2 mux_inst_3032 (
  .O(mux_o_3032),
  .I0(mux_o_3015),
  .I1(mux_o_3016),
  .S0(dff_q_4)
);
MUX2 mux_inst_3033 (
  .O(mux_o_3033),
  .I0(mux_o_3017),
  .I1(mux_o_3018),
  .S0(dff_q_3)
);
MUX2 mux_inst_3034 (
  .O(mux_o_3034),
  .I0(mux_o_3019),
  .I1(mux_o_3020),
  .S0(dff_q_3)
);
MUX2 mux_inst_3035 (
  .O(mux_o_3035),
  .I0(mux_o_3021),
  .I1(mux_o_3022),
  .S0(dff_q_3)
);
MUX2 mux_inst_3036 (
  .O(mux_o_3036),
  .I0(mux_o_3023),
  .I1(mux_o_3024),
  .S0(dff_q_3)
);
MUX2 mux_inst_3037 (
  .O(mux_o_3037),
  .I0(mux_o_3025),
  .I1(mux_o_3026),
  .S0(dff_q_3)
);
MUX2 mux_inst_3038 (
  .O(mux_o_3038),
  .I0(mux_o_3027),
  .I1(mux_o_3028),
  .S0(dff_q_3)
);
MUX2 mux_inst_3039 (
  .O(mux_o_3039),
  .I0(mux_o_3029),
  .I1(mux_o_3030),
  .S0(dff_q_3)
);
MUX2 mux_inst_3040 (
  .O(mux_o_3040),
  .I0(mux_o_3031),
  .I1(mux_o_3032),
  .S0(dff_q_3)
);
MUX2 mux_inst_3041 (
  .O(mux_o_3041),
  .I0(mux_o_3033),
  .I1(mux_o_3034),
  .S0(dff_q_2)
);
MUX2 mux_inst_3042 (
  .O(mux_o_3042),
  .I0(mux_o_3035),
  .I1(mux_o_3036),
  .S0(dff_q_2)
);
MUX2 mux_inst_3043 (
  .O(mux_o_3043),
  .I0(mux_o_3037),
  .I1(mux_o_3038),
  .S0(dff_q_2)
);
MUX2 mux_inst_3044 (
  .O(mux_o_3044),
  .I0(mux_o_3039),
  .I1(mux_o_3040),
  .S0(dff_q_2)
);
MUX2 mux_inst_3045 (
  .O(mux_o_3045),
  .I0(mux_o_3041),
  .I1(mux_o_3042),
  .S0(dff_q_1)
);
MUX2 mux_inst_3046 (
  .O(mux_o_3046),
  .I0(mux_o_3043),
  .I1(mux_o_3044),
  .S0(dff_q_1)
);
MUX2 mux_inst_3047 (
  .O(dout[23]),
  .I0(mux_o_3045),
  .I1(mux_o_3046),
  .S0(dff_q_0)
);
MUX2 mux_inst_3048 (
  .O(mux_o_3048),
  .I0(sdpb_inst_128_dout[24]),
  .I1(sdpb_inst_129_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3049 (
  .O(mux_o_3049),
  .I0(sdpb_inst_130_dout[24]),
  .I1(sdpb_inst_131_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3050 (
  .O(mux_o_3050),
  .I0(sdpb_inst_132_dout[24]),
  .I1(sdpb_inst_133_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3051 (
  .O(mux_o_3051),
  .I0(sdpb_inst_134_dout[24]),
  .I1(sdpb_inst_135_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3052 (
  .O(mux_o_3052),
  .I0(sdpb_inst_136_dout[24]),
  .I1(sdpb_inst_137_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3053 (
  .O(mux_o_3053),
  .I0(sdpb_inst_138_dout[24]),
  .I1(sdpb_inst_139_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3054 (
  .O(mux_o_3054),
  .I0(sdpb_inst_140_dout[24]),
  .I1(sdpb_inst_141_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3055 (
  .O(mux_o_3055),
  .I0(sdpb_inst_142_dout[24]),
  .I1(sdpb_inst_143_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3056 (
  .O(mux_o_3056),
  .I0(sdpb_inst_144_dout[24]),
  .I1(sdpb_inst_145_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3057 (
  .O(mux_o_3057),
  .I0(sdpb_inst_146_dout[24]),
  .I1(sdpb_inst_147_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3058 (
  .O(mux_o_3058),
  .I0(sdpb_inst_148_dout[24]),
  .I1(sdpb_inst_149_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3059 (
  .O(mux_o_3059),
  .I0(sdpb_inst_150_dout[24]),
  .I1(sdpb_inst_151_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3060 (
  .O(mux_o_3060),
  .I0(sdpb_inst_152_dout[24]),
  .I1(sdpb_inst_153_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3061 (
  .O(mux_o_3061),
  .I0(sdpb_inst_154_dout[24]),
  .I1(sdpb_inst_155_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3062 (
  .O(mux_o_3062),
  .I0(sdpb_inst_156_dout[24]),
  .I1(sdpb_inst_157_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3063 (
  .O(mux_o_3063),
  .I0(sdpb_inst_158_dout[24]),
  .I1(sdpb_inst_159_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3064 (
  .O(mux_o_3064),
  .I0(sdpb_inst_160_dout[24]),
  .I1(sdpb_inst_161_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3065 (
  .O(mux_o_3065),
  .I0(sdpb_inst_162_dout[24]),
  .I1(sdpb_inst_163_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3066 (
  .O(mux_o_3066),
  .I0(sdpb_inst_164_dout[24]),
  .I1(sdpb_inst_165_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3067 (
  .O(mux_o_3067),
  .I0(sdpb_inst_166_dout[24]),
  .I1(sdpb_inst_167_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3068 (
  .O(mux_o_3068),
  .I0(sdpb_inst_168_dout[24]),
  .I1(sdpb_inst_169_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3069 (
  .O(mux_o_3069),
  .I0(sdpb_inst_170_dout[24]),
  .I1(sdpb_inst_171_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3070 (
  .O(mux_o_3070),
  .I0(sdpb_inst_172_dout[24]),
  .I1(sdpb_inst_173_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3071 (
  .O(mux_o_3071),
  .I0(sdpb_inst_174_dout[24]),
  .I1(sdpb_inst_175_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3072 (
  .O(mux_o_3072),
  .I0(sdpb_inst_176_dout[24]),
  .I1(sdpb_inst_177_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3073 (
  .O(mux_o_3073),
  .I0(sdpb_inst_178_dout[24]),
  .I1(sdpb_inst_179_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3074 (
  .O(mux_o_3074),
  .I0(sdpb_inst_180_dout[24]),
  .I1(sdpb_inst_181_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3075 (
  .O(mux_o_3075),
  .I0(sdpb_inst_182_dout[24]),
  .I1(sdpb_inst_183_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3076 (
  .O(mux_o_3076),
  .I0(sdpb_inst_184_dout[24]),
  .I1(sdpb_inst_185_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3077 (
  .O(mux_o_3077),
  .I0(sdpb_inst_186_dout[24]),
  .I1(sdpb_inst_187_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3078 (
  .O(mux_o_3078),
  .I0(sdpb_inst_188_dout[24]),
  .I1(sdpb_inst_189_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3079 (
  .O(mux_o_3079),
  .I0(sdpb_inst_190_dout[24]),
  .I1(sdpb_inst_191_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3080 (
  .O(mux_o_3080),
  .I0(sdpb_inst_192_dout[24]),
  .I1(sdpb_inst_193_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3081 (
  .O(mux_o_3081),
  .I0(sdpb_inst_194_dout[24]),
  .I1(sdpb_inst_195_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3082 (
  .O(mux_o_3082),
  .I0(sdpb_inst_196_dout[24]),
  .I1(sdpb_inst_197_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3083 (
  .O(mux_o_3083),
  .I0(sdpb_inst_198_dout[24]),
  .I1(sdpb_inst_199_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3084 (
  .O(mux_o_3084),
  .I0(sdpb_inst_200_dout[24]),
  .I1(sdpb_inst_201_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3085 (
  .O(mux_o_3085),
  .I0(sdpb_inst_202_dout[24]),
  .I1(sdpb_inst_203_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3086 (
  .O(mux_o_3086),
  .I0(sdpb_inst_204_dout[24]),
  .I1(sdpb_inst_205_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3087 (
  .O(mux_o_3087),
  .I0(sdpb_inst_206_dout[24]),
  .I1(sdpb_inst_207_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3088 (
  .O(mux_o_3088),
  .I0(sdpb_inst_208_dout[24]),
  .I1(sdpb_inst_209_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3089 (
  .O(mux_o_3089),
  .I0(sdpb_inst_210_dout[24]),
  .I1(sdpb_inst_211_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3090 (
  .O(mux_o_3090),
  .I0(sdpb_inst_212_dout[24]),
  .I1(sdpb_inst_213_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3091 (
  .O(mux_o_3091),
  .I0(sdpb_inst_214_dout[24]),
  .I1(sdpb_inst_215_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3092 (
  .O(mux_o_3092),
  .I0(sdpb_inst_216_dout[24]),
  .I1(sdpb_inst_217_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3093 (
  .O(mux_o_3093),
  .I0(sdpb_inst_218_dout[24]),
  .I1(sdpb_inst_219_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3094 (
  .O(mux_o_3094),
  .I0(sdpb_inst_220_dout[24]),
  .I1(sdpb_inst_221_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3095 (
  .O(mux_o_3095),
  .I0(sdpb_inst_222_dout[24]),
  .I1(sdpb_inst_223_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3096 (
  .O(mux_o_3096),
  .I0(sdpb_inst_224_dout[24]),
  .I1(sdpb_inst_225_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3097 (
  .O(mux_o_3097),
  .I0(sdpb_inst_226_dout[24]),
  .I1(sdpb_inst_227_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3098 (
  .O(mux_o_3098),
  .I0(sdpb_inst_228_dout[24]),
  .I1(sdpb_inst_229_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3099 (
  .O(mux_o_3099),
  .I0(sdpb_inst_230_dout[24]),
  .I1(sdpb_inst_231_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3100 (
  .O(mux_o_3100),
  .I0(sdpb_inst_232_dout[24]),
  .I1(sdpb_inst_233_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3101 (
  .O(mux_o_3101),
  .I0(sdpb_inst_234_dout[24]),
  .I1(sdpb_inst_235_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3102 (
  .O(mux_o_3102),
  .I0(sdpb_inst_236_dout[24]),
  .I1(sdpb_inst_237_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3103 (
  .O(mux_o_3103),
  .I0(sdpb_inst_238_dout[24]),
  .I1(sdpb_inst_239_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3104 (
  .O(mux_o_3104),
  .I0(sdpb_inst_240_dout[24]),
  .I1(sdpb_inst_241_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3105 (
  .O(mux_o_3105),
  .I0(sdpb_inst_242_dout[24]),
  .I1(sdpb_inst_243_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3106 (
  .O(mux_o_3106),
  .I0(sdpb_inst_244_dout[24]),
  .I1(sdpb_inst_245_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3107 (
  .O(mux_o_3107),
  .I0(sdpb_inst_246_dout[24]),
  .I1(sdpb_inst_247_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3108 (
  .O(mux_o_3108),
  .I0(sdpb_inst_248_dout[24]),
  .I1(sdpb_inst_249_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3109 (
  .O(mux_o_3109),
  .I0(sdpb_inst_250_dout[24]),
  .I1(sdpb_inst_251_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3110 (
  .O(mux_o_3110),
  .I0(sdpb_inst_252_dout[24]),
  .I1(sdpb_inst_253_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3111 (
  .O(mux_o_3111),
  .I0(sdpb_inst_254_dout[24]),
  .I1(sdpb_inst_255_dout[24]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3112 (
  .O(mux_o_3112),
  .I0(mux_o_3048),
  .I1(mux_o_3049),
  .S0(dff_q_5)
);
MUX2 mux_inst_3113 (
  .O(mux_o_3113),
  .I0(mux_o_3050),
  .I1(mux_o_3051),
  .S0(dff_q_5)
);
MUX2 mux_inst_3114 (
  .O(mux_o_3114),
  .I0(mux_o_3052),
  .I1(mux_o_3053),
  .S0(dff_q_5)
);
MUX2 mux_inst_3115 (
  .O(mux_o_3115),
  .I0(mux_o_3054),
  .I1(mux_o_3055),
  .S0(dff_q_5)
);
MUX2 mux_inst_3116 (
  .O(mux_o_3116),
  .I0(mux_o_3056),
  .I1(mux_o_3057),
  .S0(dff_q_5)
);
MUX2 mux_inst_3117 (
  .O(mux_o_3117),
  .I0(mux_o_3058),
  .I1(mux_o_3059),
  .S0(dff_q_5)
);
MUX2 mux_inst_3118 (
  .O(mux_o_3118),
  .I0(mux_o_3060),
  .I1(mux_o_3061),
  .S0(dff_q_5)
);
MUX2 mux_inst_3119 (
  .O(mux_o_3119),
  .I0(mux_o_3062),
  .I1(mux_o_3063),
  .S0(dff_q_5)
);
MUX2 mux_inst_3120 (
  .O(mux_o_3120),
  .I0(mux_o_3064),
  .I1(mux_o_3065),
  .S0(dff_q_5)
);
MUX2 mux_inst_3121 (
  .O(mux_o_3121),
  .I0(mux_o_3066),
  .I1(mux_o_3067),
  .S0(dff_q_5)
);
MUX2 mux_inst_3122 (
  .O(mux_o_3122),
  .I0(mux_o_3068),
  .I1(mux_o_3069),
  .S0(dff_q_5)
);
MUX2 mux_inst_3123 (
  .O(mux_o_3123),
  .I0(mux_o_3070),
  .I1(mux_o_3071),
  .S0(dff_q_5)
);
MUX2 mux_inst_3124 (
  .O(mux_o_3124),
  .I0(mux_o_3072),
  .I1(mux_o_3073),
  .S0(dff_q_5)
);
MUX2 mux_inst_3125 (
  .O(mux_o_3125),
  .I0(mux_o_3074),
  .I1(mux_o_3075),
  .S0(dff_q_5)
);
MUX2 mux_inst_3126 (
  .O(mux_o_3126),
  .I0(mux_o_3076),
  .I1(mux_o_3077),
  .S0(dff_q_5)
);
MUX2 mux_inst_3127 (
  .O(mux_o_3127),
  .I0(mux_o_3078),
  .I1(mux_o_3079),
  .S0(dff_q_5)
);
MUX2 mux_inst_3128 (
  .O(mux_o_3128),
  .I0(mux_o_3080),
  .I1(mux_o_3081),
  .S0(dff_q_5)
);
MUX2 mux_inst_3129 (
  .O(mux_o_3129),
  .I0(mux_o_3082),
  .I1(mux_o_3083),
  .S0(dff_q_5)
);
MUX2 mux_inst_3130 (
  .O(mux_o_3130),
  .I0(mux_o_3084),
  .I1(mux_o_3085),
  .S0(dff_q_5)
);
MUX2 mux_inst_3131 (
  .O(mux_o_3131),
  .I0(mux_o_3086),
  .I1(mux_o_3087),
  .S0(dff_q_5)
);
MUX2 mux_inst_3132 (
  .O(mux_o_3132),
  .I0(mux_o_3088),
  .I1(mux_o_3089),
  .S0(dff_q_5)
);
MUX2 mux_inst_3133 (
  .O(mux_o_3133),
  .I0(mux_o_3090),
  .I1(mux_o_3091),
  .S0(dff_q_5)
);
MUX2 mux_inst_3134 (
  .O(mux_o_3134),
  .I0(mux_o_3092),
  .I1(mux_o_3093),
  .S0(dff_q_5)
);
MUX2 mux_inst_3135 (
  .O(mux_o_3135),
  .I0(mux_o_3094),
  .I1(mux_o_3095),
  .S0(dff_q_5)
);
MUX2 mux_inst_3136 (
  .O(mux_o_3136),
  .I0(mux_o_3096),
  .I1(mux_o_3097),
  .S0(dff_q_5)
);
MUX2 mux_inst_3137 (
  .O(mux_o_3137),
  .I0(mux_o_3098),
  .I1(mux_o_3099),
  .S0(dff_q_5)
);
MUX2 mux_inst_3138 (
  .O(mux_o_3138),
  .I0(mux_o_3100),
  .I1(mux_o_3101),
  .S0(dff_q_5)
);
MUX2 mux_inst_3139 (
  .O(mux_o_3139),
  .I0(mux_o_3102),
  .I1(mux_o_3103),
  .S0(dff_q_5)
);
MUX2 mux_inst_3140 (
  .O(mux_o_3140),
  .I0(mux_o_3104),
  .I1(mux_o_3105),
  .S0(dff_q_5)
);
MUX2 mux_inst_3141 (
  .O(mux_o_3141),
  .I0(mux_o_3106),
  .I1(mux_o_3107),
  .S0(dff_q_5)
);
MUX2 mux_inst_3142 (
  .O(mux_o_3142),
  .I0(mux_o_3108),
  .I1(mux_o_3109),
  .S0(dff_q_5)
);
MUX2 mux_inst_3143 (
  .O(mux_o_3143),
  .I0(mux_o_3110),
  .I1(mux_o_3111),
  .S0(dff_q_5)
);
MUX2 mux_inst_3144 (
  .O(mux_o_3144),
  .I0(mux_o_3112),
  .I1(mux_o_3113),
  .S0(dff_q_4)
);
MUX2 mux_inst_3145 (
  .O(mux_o_3145),
  .I0(mux_o_3114),
  .I1(mux_o_3115),
  .S0(dff_q_4)
);
MUX2 mux_inst_3146 (
  .O(mux_o_3146),
  .I0(mux_o_3116),
  .I1(mux_o_3117),
  .S0(dff_q_4)
);
MUX2 mux_inst_3147 (
  .O(mux_o_3147),
  .I0(mux_o_3118),
  .I1(mux_o_3119),
  .S0(dff_q_4)
);
MUX2 mux_inst_3148 (
  .O(mux_o_3148),
  .I0(mux_o_3120),
  .I1(mux_o_3121),
  .S0(dff_q_4)
);
MUX2 mux_inst_3149 (
  .O(mux_o_3149),
  .I0(mux_o_3122),
  .I1(mux_o_3123),
  .S0(dff_q_4)
);
MUX2 mux_inst_3150 (
  .O(mux_o_3150),
  .I0(mux_o_3124),
  .I1(mux_o_3125),
  .S0(dff_q_4)
);
MUX2 mux_inst_3151 (
  .O(mux_o_3151),
  .I0(mux_o_3126),
  .I1(mux_o_3127),
  .S0(dff_q_4)
);
MUX2 mux_inst_3152 (
  .O(mux_o_3152),
  .I0(mux_o_3128),
  .I1(mux_o_3129),
  .S0(dff_q_4)
);
MUX2 mux_inst_3153 (
  .O(mux_o_3153),
  .I0(mux_o_3130),
  .I1(mux_o_3131),
  .S0(dff_q_4)
);
MUX2 mux_inst_3154 (
  .O(mux_o_3154),
  .I0(mux_o_3132),
  .I1(mux_o_3133),
  .S0(dff_q_4)
);
MUX2 mux_inst_3155 (
  .O(mux_o_3155),
  .I0(mux_o_3134),
  .I1(mux_o_3135),
  .S0(dff_q_4)
);
MUX2 mux_inst_3156 (
  .O(mux_o_3156),
  .I0(mux_o_3136),
  .I1(mux_o_3137),
  .S0(dff_q_4)
);
MUX2 mux_inst_3157 (
  .O(mux_o_3157),
  .I0(mux_o_3138),
  .I1(mux_o_3139),
  .S0(dff_q_4)
);
MUX2 mux_inst_3158 (
  .O(mux_o_3158),
  .I0(mux_o_3140),
  .I1(mux_o_3141),
  .S0(dff_q_4)
);
MUX2 mux_inst_3159 (
  .O(mux_o_3159),
  .I0(mux_o_3142),
  .I1(mux_o_3143),
  .S0(dff_q_4)
);
MUX2 mux_inst_3160 (
  .O(mux_o_3160),
  .I0(mux_o_3144),
  .I1(mux_o_3145),
  .S0(dff_q_3)
);
MUX2 mux_inst_3161 (
  .O(mux_o_3161),
  .I0(mux_o_3146),
  .I1(mux_o_3147),
  .S0(dff_q_3)
);
MUX2 mux_inst_3162 (
  .O(mux_o_3162),
  .I0(mux_o_3148),
  .I1(mux_o_3149),
  .S0(dff_q_3)
);
MUX2 mux_inst_3163 (
  .O(mux_o_3163),
  .I0(mux_o_3150),
  .I1(mux_o_3151),
  .S0(dff_q_3)
);
MUX2 mux_inst_3164 (
  .O(mux_o_3164),
  .I0(mux_o_3152),
  .I1(mux_o_3153),
  .S0(dff_q_3)
);
MUX2 mux_inst_3165 (
  .O(mux_o_3165),
  .I0(mux_o_3154),
  .I1(mux_o_3155),
  .S0(dff_q_3)
);
MUX2 mux_inst_3166 (
  .O(mux_o_3166),
  .I0(mux_o_3156),
  .I1(mux_o_3157),
  .S0(dff_q_3)
);
MUX2 mux_inst_3167 (
  .O(mux_o_3167),
  .I0(mux_o_3158),
  .I1(mux_o_3159),
  .S0(dff_q_3)
);
MUX2 mux_inst_3168 (
  .O(mux_o_3168),
  .I0(mux_o_3160),
  .I1(mux_o_3161),
  .S0(dff_q_2)
);
MUX2 mux_inst_3169 (
  .O(mux_o_3169),
  .I0(mux_o_3162),
  .I1(mux_o_3163),
  .S0(dff_q_2)
);
MUX2 mux_inst_3170 (
  .O(mux_o_3170),
  .I0(mux_o_3164),
  .I1(mux_o_3165),
  .S0(dff_q_2)
);
MUX2 mux_inst_3171 (
  .O(mux_o_3171),
  .I0(mux_o_3166),
  .I1(mux_o_3167),
  .S0(dff_q_2)
);
MUX2 mux_inst_3172 (
  .O(mux_o_3172),
  .I0(mux_o_3168),
  .I1(mux_o_3169),
  .S0(dff_q_1)
);
MUX2 mux_inst_3173 (
  .O(mux_o_3173),
  .I0(mux_o_3170),
  .I1(mux_o_3171),
  .S0(dff_q_1)
);
MUX2 mux_inst_3174 (
  .O(dout[24]),
  .I0(mux_o_3172),
  .I1(mux_o_3173),
  .S0(dff_q_0)
);
MUX2 mux_inst_3175 (
  .O(mux_o_3175),
  .I0(sdpb_inst_128_dout[25]),
  .I1(sdpb_inst_129_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3176 (
  .O(mux_o_3176),
  .I0(sdpb_inst_130_dout[25]),
  .I1(sdpb_inst_131_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3177 (
  .O(mux_o_3177),
  .I0(sdpb_inst_132_dout[25]),
  .I1(sdpb_inst_133_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3178 (
  .O(mux_o_3178),
  .I0(sdpb_inst_134_dout[25]),
  .I1(sdpb_inst_135_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3179 (
  .O(mux_o_3179),
  .I0(sdpb_inst_136_dout[25]),
  .I1(sdpb_inst_137_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3180 (
  .O(mux_o_3180),
  .I0(sdpb_inst_138_dout[25]),
  .I1(sdpb_inst_139_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3181 (
  .O(mux_o_3181),
  .I0(sdpb_inst_140_dout[25]),
  .I1(sdpb_inst_141_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3182 (
  .O(mux_o_3182),
  .I0(sdpb_inst_142_dout[25]),
  .I1(sdpb_inst_143_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3183 (
  .O(mux_o_3183),
  .I0(sdpb_inst_144_dout[25]),
  .I1(sdpb_inst_145_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3184 (
  .O(mux_o_3184),
  .I0(sdpb_inst_146_dout[25]),
  .I1(sdpb_inst_147_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3185 (
  .O(mux_o_3185),
  .I0(sdpb_inst_148_dout[25]),
  .I1(sdpb_inst_149_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3186 (
  .O(mux_o_3186),
  .I0(sdpb_inst_150_dout[25]),
  .I1(sdpb_inst_151_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3187 (
  .O(mux_o_3187),
  .I0(sdpb_inst_152_dout[25]),
  .I1(sdpb_inst_153_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3188 (
  .O(mux_o_3188),
  .I0(sdpb_inst_154_dout[25]),
  .I1(sdpb_inst_155_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3189 (
  .O(mux_o_3189),
  .I0(sdpb_inst_156_dout[25]),
  .I1(sdpb_inst_157_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3190 (
  .O(mux_o_3190),
  .I0(sdpb_inst_158_dout[25]),
  .I1(sdpb_inst_159_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3191 (
  .O(mux_o_3191),
  .I0(sdpb_inst_160_dout[25]),
  .I1(sdpb_inst_161_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3192 (
  .O(mux_o_3192),
  .I0(sdpb_inst_162_dout[25]),
  .I1(sdpb_inst_163_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3193 (
  .O(mux_o_3193),
  .I0(sdpb_inst_164_dout[25]),
  .I1(sdpb_inst_165_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3194 (
  .O(mux_o_3194),
  .I0(sdpb_inst_166_dout[25]),
  .I1(sdpb_inst_167_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3195 (
  .O(mux_o_3195),
  .I0(sdpb_inst_168_dout[25]),
  .I1(sdpb_inst_169_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3196 (
  .O(mux_o_3196),
  .I0(sdpb_inst_170_dout[25]),
  .I1(sdpb_inst_171_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3197 (
  .O(mux_o_3197),
  .I0(sdpb_inst_172_dout[25]),
  .I1(sdpb_inst_173_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3198 (
  .O(mux_o_3198),
  .I0(sdpb_inst_174_dout[25]),
  .I1(sdpb_inst_175_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3199 (
  .O(mux_o_3199),
  .I0(sdpb_inst_176_dout[25]),
  .I1(sdpb_inst_177_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3200 (
  .O(mux_o_3200),
  .I0(sdpb_inst_178_dout[25]),
  .I1(sdpb_inst_179_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3201 (
  .O(mux_o_3201),
  .I0(sdpb_inst_180_dout[25]),
  .I1(sdpb_inst_181_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3202 (
  .O(mux_o_3202),
  .I0(sdpb_inst_182_dout[25]),
  .I1(sdpb_inst_183_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3203 (
  .O(mux_o_3203),
  .I0(sdpb_inst_184_dout[25]),
  .I1(sdpb_inst_185_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3204 (
  .O(mux_o_3204),
  .I0(sdpb_inst_186_dout[25]),
  .I1(sdpb_inst_187_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3205 (
  .O(mux_o_3205),
  .I0(sdpb_inst_188_dout[25]),
  .I1(sdpb_inst_189_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3206 (
  .O(mux_o_3206),
  .I0(sdpb_inst_190_dout[25]),
  .I1(sdpb_inst_191_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3207 (
  .O(mux_o_3207),
  .I0(sdpb_inst_192_dout[25]),
  .I1(sdpb_inst_193_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3208 (
  .O(mux_o_3208),
  .I0(sdpb_inst_194_dout[25]),
  .I1(sdpb_inst_195_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3209 (
  .O(mux_o_3209),
  .I0(sdpb_inst_196_dout[25]),
  .I1(sdpb_inst_197_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3210 (
  .O(mux_o_3210),
  .I0(sdpb_inst_198_dout[25]),
  .I1(sdpb_inst_199_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3211 (
  .O(mux_o_3211),
  .I0(sdpb_inst_200_dout[25]),
  .I1(sdpb_inst_201_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3212 (
  .O(mux_o_3212),
  .I0(sdpb_inst_202_dout[25]),
  .I1(sdpb_inst_203_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3213 (
  .O(mux_o_3213),
  .I0(sdpb_inst_204_dout[25]),
  .I1(sdpb_inst_205_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3214 (
  .O(mux_o_3214),
  .I0(sdpb_inst_206_dout[25]),
  .I1(sdpb_inst_207_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3215 (
  .O(mux_o_3215),
  .I0(sdpb_inst_208_dout[25]),
  .I1(sdpb_inst_209_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3216 (
  .O(mux_o_3216),
  .I0(sdpb_inst_210_dout[25]),
  .I1(sdpb_inst_211_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3217 (
  .O(mux_o_3217),
  .I0(sdpb_inst_212_dout[25]),
  .I1(sdpb_inst_213_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3218 (
  .O(mux_o_3218),
  .I0(sdpb_inst_214_dout[25]),
  .I1(sdpb_inst_215_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3219 (
  .O(mux_o_3219),
  .I0(sdpb_inst_216_dout[25]),
  .I1(sdpb_inst_217_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3220 (
  .O(mux_o_3220),
  .I0(sdpb_inst_218_dout[25]),
  .I1(sdpb_inst_219_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3221 (
  .O(mux_o_3221),
  .I0(sdpb_inst_220_dout[25]),
  .I1(sdpb_inst_221_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3222 (
  .O(mux_o_3222),
  .I0(sdpb_inst_222_dout[25]),
  .I1(sdpb_inst_223_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3223 (
  .O(mux_o_3223),
  .I0(sdpb_inst_224_dout[25]),
  .I1(sdpb_inst_225_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3224 (
  .O(mux_o_3224),
  .I0(sdpb_inst_226_dout[25]),
  .I1(sdpb_inst_227_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3225 (
  .O(mux_o_3225),
  .I0(sdpb_inst_228_dout[25]),
  .I1(sdpb_inst_229_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3226 (
  .O(mux_o_3226),
  .I0(sdpb_inst_230_dout[25]),
  .I1(sdpb_inst_231_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3227 (
  .O(mux_o_3227),
  .I0(sdpb_inst_232_dout[25]),
  .I1(sdpb_inst_233_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3228 (
  .O(mux_o_3228),
  .I0(sdpb_inst_234_dout[25]),
  .I1(sdpb_inst_235_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3229 (
  .O(mux_o_3229),
  .I0(sdpb_inst_236_dout[25]),
  .I1(sdpb_inst_237_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3230 (
  .O(mux_o_3230),
  .I0(sdpb_inst_238_dout[25]),
  .I1(sdpb_inst_239_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3231 (
  .O(mux_o_3231),
  .I0(sdpb_inst_240_dout[25]),
  .I1(sdpb_inst_241_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3232 (
  .O(mux_o_3232),
  .I0(sdpb_inst_242_dout[25]),
  .I1(sdpb_inst_243_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3233 (
  .O(mux_o_3233),
  .I0(sdpb_inst_244_dout[25]),
  .I1(sdpb_inst_245_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3234 (
  .O(mux_o_3234),
  .I0(sdpb_inst_246_dout[25]),
  .I1(sdpb_inst_247_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3235 (
  .O(mux_o_3235),
  .I0(sdpb_inst_248_dout[25]),
  .I1(sdpb_inst_249_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3236 (
  .O(mux_o_3236),
  .I0(sdpb_inst_250_dout[25]),
  .I1(sdpb_inst_251_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3237 (
  .O(mux_o_3237),
  .I0(sdpb_inst_252_dout[25]),
  .I1(sdpb_inst_253_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3238 (
  .O(mux_o_3238),
  .I0(sdpb_inst_254_dout[25]),
  .I1(sdpb_inst_255_dout[25]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3239 (
  .O(mux_o_3239),
  .I0(mux_o_3175),
  .I1(mux_o_3176),
  .S0(dff_q_5)
);
MUX2 mux_inst_3240 (
  .O(mux_o_3240),
  .I0(mux_o_3177),
  .I1(mux_o_3178),
  .S0(dff_q_5)
);
MUX2 mux_inst_3241 (
  .O(mux_o_3241),
  .I0(mux_o_3179),
  .I1(mux_o_3180),
  .S0(dff_q_5)
);
MUX2 mux_inst_3242 (
  .O(mux_o_3242),
  .I0(mux_o_3181),
  .I1(mux_o_3182),
  .S0(dff_q_5)
);
MUX2 mux_inst_3243 (
  .O(mux_o_3243),
  .I0(mux_o_3183),
  .I1(mux_o_3184),
  .S0(dff_q_5)
);
MUX2 mux_inst_3244 (
  .O(mux_o_3244),
  .I0(mux_o_3185),
  .I1(mux_o_3186),
  .S0(dff_q_5)
);
MUX2 mux_inst_3245 (
  .O(mux_o_3245),
  .I0(mux_o_3187),
  .I1(mux_o_3188),
  .S0(dff_q_5)
);
MUX2 mux_inst_3246 (
  .O(mux_o_3246),
  .I0(mux_o_3189),
  .I1(mux_o_3190),
  .S0(dff_q_5)
);
MUX2 mux_inst_3247 (
  .O(mux_o_3247),
  .I0(mux_o_3191),
  .I1(mux_o_3192),
  .S0(dff_q_5)
);
MUX2 mux_inst_3248 (
  .O(mux_o_3248),
  .I0(mux_o_3193),
  .I1(mux_o_3194),
  .S0(dff_q_5)
);
MUX2 mux_inst_3249 (
  .O(mux_o_3249),
  .I0(mux_o_3195),
  .I1(mux_o_3196),
  .S0(dff_q_5)
);
MUX2 mux_inst_3250 (
  .O(mux_o_3250),
  .I0(mux_o_3197),
  .I1(mux_o_3198),
  .S0(dff_q_5)
);
MUX2 mux_inst_3251 (
  .O(mux_o_3251),
  .I0(mux_o_3199),
  .I1(mux_o_3200),
  .S0(dff_q_5)
);
MUX2 mux_inst_3252 (
  .O(mux_o_3252),
  .I0(mux_o_3201),
  .I1(mux_o_3202),
  .S0(dff_q_5)
);
MUX2 mux_inst_3253 (
  .O(mux_o_3253),
  .I0(mux_o_3203),
  .I1(mux_o_3204),
  .S0(dff_q_5)
);
MUX2 mux_inst_3254 (
  .O(mux_o_3254),
  .I0(mux_o_3205),
  .I1(mux_o_3206),
  .S0(dff_q_5)
);
MUX2 mux_inst_3255 (
  .O(mux_o_3255),
  .I0(mux_o_3207),
  .I1(mux_o_3208),
  .S0(dff_q_5)
);
MUX2 mux_inst_3256 (
  .O(mux_o_3256),
  .I0(mux_o_3209),
  .I1(mux_o_3210),
  .S0(dff_q_5)
);
MUX2 mux_inst_3257 (
  .O(mux_o_3257),
  .I0(mux_o_3211),
  .I1(mux_o_3212),
  .S0(dff_q_5)
);
MUX2 mux_inst_3258 (
  .O(mux_o_3258),
  .I0(mux_o_3213),
  .I1(mux_o_3214),
  .S0(dff_q_5)
);
MUX2 mux_inst_3259 (
  .O(mux_o_3259),
  .I0(mux_o_3215),
  .I1(mux_o_3216),
  .S0(dff_q_5)
);
MUX2 mux_inst_3260 (
  .O(mux_o_3260),
  .I0(mux_o_3217),
  .I1(mux_o_3218),
  .S0(dff_q_5)
);
MUX2 mux_inst_3261 (
  .O(mux_o_3261),
  .I0(mux_o_3219),
  .I1(mux_o_3220),
  .S0(dff_q_5)
);
MUX2 mux_inst_3262 (
  .O(mux_o_3262),
  .I0(mux_o_3221),
  .I1(mux_o_3222),
  .S0(dff_q_5)
);
MUX2 mux_inst_3263 (
  .O(mux_o_3263),
  .I0(mux_o_3223),
  .I1(mux_o_3224),
  .S0(dff_q_5)
);
MUX2 mux_inst_3264 (
  .O(mux_o_3264),
  .I0(mux_o_3225),
  .I1(mux_o_3226),
  .S0(dff_q_5)
);
MUX2 mux_inst_3265 (
  .O(mux_o_3265),
  .I0(mux_o_3227),
  .I1(mux_o_3228),
  .S0(dff_q_5)
);
MUX2 mux_inst_3266 (
  .O(mux_o_3266),
  .I0(mux_o_3229),
  .I1(mux_o_3230),
  .S0(dff_q_5)
);
MUX2 mux_inst_3267 (
  .O(mux_o_3267),
  .I0(mux_o_3231),
  .I1(mux_o_3232),
  .S0(dff_q_5)
);
MUX2 mux_inst_3268 (
  .O(mux_o_3268),
  .I0(mux_o_3233),
  .I1(mux_o_3234),
  .S0(dff_q_5)
);
MUX2 mux_inst_3269 (
  .O(mux_o_3269),
  .I0(mux_o_3235),
  .I1(mux_o_3236),
  .S0(dff_q_5)
);
MUX2 mux_inst_3270 (
  .O(mux_o_3270),
  .I0(mux_o_3237),
  .I1(mux_o_3238),
  .S0(dff_q_5)
);
MUX2 mux_inst_3271 (
  .O(mux_o_3271),
  .I0(mux_o_3239),
  .I1(mux_o_3240),
  .S0(dff_q_4)
);
MUX2 mux_inst_3272 (
  .O(mux_o_3272),
  .I0(mux_o_3241),
  .I1(mux_o_3242),
  .S0(dff_q_4)
);
MUX2 mux_inst_3273 (
  .O(mux_o_3273),
  .I0(mux_o_3243),
  .I1(mux_o_3244),
  .S0(dff_q_4)
);
MUX2 mux_inst_3274 (
  .O(mux_o_3274),
  .I0(mux_o_3245),
  .I1(mux_o_3246),
  .S0(dff_q_4)
);
MUX2 mux_inst_3275 (
  .O(mux_o_3275),
  .I0(mux_o_3247),
  .I1(mux_o_3248),
  .S0(dff_q_4)
);
MUX2 mux_inst_3276 (
  .O(mux_o_3276),
  .I0(mux_o_3249),
  .I1(mux_o_3250),
  .S0(dff_q_4)
);
MUX2 mux_inst_3277 (
  .O(mux_o_3277),
  .I0(mux_o_3251),
  .I1(mux_o_3252),
  .S0(dff_q_4)
);
MUX2 mux_inst_3278 (
  .O(mux_o_3278),
  .I0(mux_o_3253),
  .I1(mux_o_3254),
  .S0(dff_q_4)
);
MUX2 mux_inst_3279 (
  .O(mux_o_3279),
  .I0(mux_o_3255),
  .I1(mux_o_3256),
  .S0(dff_q_4)
);
MUX2 mux_inst_3280 (
  .O(mux_o_3280),
  .I0(mux_o_3257),
  .I1(mux_o_3258),
  .S0(dff_q_4)
);
MUX2 mux_inst_3281 (
  .O(mux_o_3281),
  .I0(mux_o_3259),
  .I1(mux_o_3260),
  .S0(dff_q_4)
);
MUX2 mux_inst_3282 (
  .O(mux_o_3282),
  .I0(mux_o_3261),
  .I1(mux_o_3262),
  .S0(dff_q_4)
);
MUX2 mux_inst_3283 (
  .O(mux_o_3283),
  .I0(mux_o_3263),
  .I1(mux_o_3264),
  .S0(dff_q_4)
);
MUX2 mux_inst_3284 (
  .O(mux_o_3284),
  .I0(mux_o_3265),
  .I1(mux_o_3266),
  .S0(dff_q_4)
);
MUX2 mux_inst_3285 (
  .O(mux_o_3285),
  .I0(mux_o_3267),
  .I1(mux_o_3268),
  .S0(dff_q_4)
);
MUX2 mux_inst_3286 (
  .O(mux_o_3286),
  .I0(mux_o_3269),
  .I1(mux_o_3270),
  .S0(dff_q_4)
);
MUX2 mux_inst_3287 (
  .O(mux_o_3287),
  .I0(mux_o_3271),
  .I1(mux_o_3272),
  .S0(dff_q_3)
);
MUX2 mux_inst_3288 (
  .O(mux_o_3288),
  .I0(mux_o_3273),
  .I1(mux_o_3274),
  .S0(dff_q_3)
);
MUX2 mux_inst_3289 (
  .O(mux_o_3289),
  .I0(mux_o_3275),
  .I1(mux_o_3276),
  .S0(dff_q_3)
);
MUX2 mux_inst_3290 (
  .O(mux_o_3290),
  .I0(mux_o_3277),
  .I1(mux_o_3278),
  .S0(dff_q_3)
);
MUX2 mux_inst_3291 (
  .O(mux_o_3291),
  .I0(mux_o_3279),
  .I1(mux_o_3280),
  .S0(dff_q_3)
);
MUX2 mux_inst_3292 (
  .O(mux_o_3292),
  .I0(mux_o_3281),
  .I1(mux_o_3282),
  .S0(dff_q_3)
);
MUX2 mux_inst_3293 (
  .O(mux_o_3293),
  .I0(mux_o_3283),
  .I1(mux_o_3284),
  .S0(dff_q_3)
);
MUX2 mux_inst_3294 (
  .O(mux_o_3294),
  .I0(mux_o_3285),
  .I1(mux_o_3286),
  .S0(dff_q_3)
);
MUX2 mux_inst_3295 (
  .O(mux_o_3295),
  .I0(mux_o_3287),
  .I1(mux_o_3288),
  .S0(dff_q_2)
);
MUX2 mux_inst_3296 (
  .O(mux_o_3296),
  .I0(mux_o_3289),
  .I1(mux_o_3290),
  .S0(dff_q_2)
);
MUX2 mux_inst_3297 (
  .O(mux_o_3297),
  .I0(mux_o_3291),
  .I1(mux_o_3292),
  .S0(dff_q_2)
);
MUX2 mux_inst_3298 (
  .O(mux_o_3298),
  .I0(mux_o_3293),
  .I1(mux_o_3294),
  .S0(dff_q_2)
);
MUX2 mux_inst_3299 (
  .O(mux_o_3299),
  .I0(mux_o_3295),
  .I1(mux_o_3296),
  .S0(dff_q_1)
);
MUX2 mux_inst_3300 (
  .O(mux_o_3300),
  .I0(mux_o_3297),
  .I1(mux_o_3298),
  .S0(dff_q_1)
);
MUX2 mux_inst_3301 (
  .O(dout[25]),
  .I0(mux_o_3299),
  .I1(mux_o_3300),
  .S0(dff_q_0)
);
MUX2 mux_inst_3302 (
  .O(mux_o_3302),
  .I0(sdpb_inst_128_dout[26]),
  .I1(sdpb_inst_129_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3303 (
  .O(mux_o_3303),
  .I0(sdpb_inst_130_dout[26]),
  .I1(sdpb_inst_131_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3304 (
  .O(mux_o_3304),
  .I0(sdpb_inst_132_dout[26]),
  .I1(sdpb_inst_133_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3305 (
  .O(mux_o_3305),
  .I0(sdpb_inst_134_dout[26]),
  .I1(sdpb_inst_135_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3306 (
  .O(mux_o_3306),
  .I0(sdpb_inst_136_dout[26]),
  .I1(sdpb_inst_137_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3307 (
  .O(mux_o_3307),
  .I0(sdpb_inst_138_dout[26]),
  .I1(sdpb_inst_139_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3308 (
  .O(mux_o_3308),
  .I0(sdpb_inst_140_dout[26]),
  .I1(sdpb_inst_141_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3309 (
  .O(mux_o_3309),
  .I0(sdpb_inst_142_dout[26]),
  .I1(sdpb_inst_143_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3310 (
  .O(mux_o_3310),
  .I0(sdpb_inst_144_dout[26]),
  .I1(sdpb_inst_145_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3311 (
  .O(mux_o_3311),
  .I0(sdpb_inst_146_dout[26]),
  .I1(sdpb_inst_147_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3312 (
  .O(mux_o_3312),
  .I0(sdpb_inst_148_dout[26]),
  .I1(sdpb_inst_149_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3313 (
  .O(mux_o_3313),
  .I0(sdpb_inst_150_dout[26]),
  .I1(sdpb_inst_151_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3314 (
  .O(mux_o_3314),
  .I0(sdpb_inst_152_dout[26]),
  .I1(sdpb_inst_153_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3315 (
  .O(mux_o_3315),
  .I0(sdpb_inst_154_dout[26]),
  .I1(sdpb_inst_155_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3316 (
  .O(mux_o_3316),
  .I0(sdpb_inst_156_dout[26]),
  .I1(sdpb_inst_157_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3317 (
  .O(mux_o_3317),
  .I0(sdpb_inst_158_dout[26]),
  .I1(sdpb_inst_159_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3318 (
  .O(mux_o_3318),
  .I0(sdpb_inst_160_dout[26]),
  .I1(sdpb_inst_161_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3319 (
  .O(mux_o_3319),
  .I0(sdpb_inst_162_dout[26]),
  .I1(sdpb_inst_163_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3320 (
  .O(mux_o_3320),
  .I0(sdpb_inst_164_dout[26]),
  .I1(sdpb_inst_165_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3321 (
  .O(mux_o_3321),
  .I0(sdpb_inst_166_dout[26]),
  .I1(sdpb_inst_167_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3322 (
  .O(mux_o_3322),
  .I0(sdpb_inst_168_dout[26]),
  .I1(sdpb_inst_169_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3323 (
  .O(mux_o_3323),
  .I0(sdpb_inst_170_dout[26]),
  .I1(sdpb_inst_171_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3324 (
  .O(mux_o_3324),
  .I0(sdpb_inst_172_dout[26]),
  .I1(sdpb_inst_173_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3325 (
  .O(mux_o_3325),
  .I0(sdpb_inst_174_dout[26]),
  .I1(sdpb_inst_175_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3326 (
  .O(mux_o_3326),
  .I0(sdpb_inst_176_dout[26]),
  .I1(sdpb_inst_177_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3327 (
  .O(mux_o_3327),
  .I0(sdpb_inst_178_dout[26]),
  .I1(sdpb_inst_179_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3328 (
  .O(mux_o_3328),
  .I0(sdpb_inst_180_dout[26]),
  .I1(sdpb_inst_181_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3329 (
  .O(mux_o_3329),
  .I0(sdpb_inst_182_dout[26]),
  .I1(sdpb_inst_183_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3330 (
  .O(mux_o_3330),
  .I0(sdpb_inst_184_dout[26]),
  .I1(sdpb_inst_185_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3331 (
  .O(mux_o_3331),
  .I0(sdpb_inst_186_dout[26]),
  .I1(sdpb_inst_187_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3332 (
  .O(mux_o_3332),
  .I0(sdpb_inst_188_dout[26]),
  .I1(sdpb_inst_189_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3333 (
  .O(mux_o_3333),
  .I0(sdpb_inst_190_dout[26]),
  .I1(sdpb_inst_191_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3334 (
  .O(mux_o_3334),
  .I0(sdpb_inst_192_dout[26]),
  .I1(sdpb_inst_193_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3335 (
  .O(mux_o_3335),
  .I0(sdpb_inst_194_dout[26]),
  .I1(sdpb_inst_195_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3336 (
  .O(mux_o_3336),
  .I0(sdpb_inst_196_dout[26]),
  .I1(sdpb_inst_197_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3337 (
  .O(mux_o_3337),
  .I0(sdpb_inst_198_dout[26]),
  .I1(sdpb_inst_199_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3338 (
  .O(mux_o_3338),
  .I0(sdpb_inst_200_dout[26]),
  .I1(sdpb_inst_201_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3339 (
  .O(mux_o_3339),
  .I0(sdpb_inst_202_dout[26]),
  .I1(sdpb_inst_203_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3340 (
  .O(mux_o_3340),
  .I0(sdpb_inst_204_dout[26]),
  .I1(sdpb_inst_205_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3341 (
  .O(mux_o_3341),
  .I0(sdpb_inst_206_dout[26]),
  .I1(sdpb_inst_207_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3342 (
  .O(mux_o_3342),
  .I0(sdpb_inst_208_dout[26]),
  .I1(sdpb_inst_209_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3343 (
  .O(mux_o_3343),
  .I0(sdpb_inst_210_dout[26]),
  .I1(sdpb_inst_211_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3344 (
  .O(mux_o_3344),
  .I0(sdpb_inst_212_dout[26]),
  .I1(sdpb_inst_213_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3345 (
  .O(mux_o_3345),
  .I0(sdpb_inst_214_dout[26]),
  .I1(sdpb_inst_215_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3346 (
  .O(mux_o_3346),
  .I0(sdpb_inst_216_dout[26]),
  .I1(sdpb_inst_217_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3347 (
  .O(mux_o_3347),
  .I0(sdpb_inst_218_dout[26]),
  .I1(sdpb_inst_219_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3348 (
  .O(mux_o_3348),
  .I0(sdpb_inst_220_dout[26]),
  .I1(sdpb_inst_221_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3349 (
  .O(mux_o_3349),
  .I0(sdpb_inst_222_dout[26]),
  .I1(sdpb_inst_223_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3350 (
  .O(mux_o_3350),
  .I0(sdpb_inst_224_dout[26]),
  .I1(sdpb_inst_225_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3351 (
  .O(mux_o_3351),
  .I0(sdpb_inst_226_dout[26]),
  .I1(sdpb_inst_227_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3352 (
  .O(mux_o_3352),
  .I0(sdpb_inst_228_dout[26]),
  .I1(sdpb_inst_229_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3353 (
  .O(mux_o_3353),
  .I0(sdpb_inst_230_dout[26]),
  .I1(sdpb_inst_231_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3354 (
  .O(mux_o_3354),
  .I0(sdpb_inst_232_dout[26]),
  .I1(sdpb_inst_233_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3355 (
  .O(mux_o_3355),
  .I0(sdpb_inst_234_dout[26]),
  .I1(sdpb_inst_235_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3356 (
  .O(mux_o_3356),
  .I0(sdpb_inst_236_dout[26]),
  .I1(sdpb_inst_237_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3357 (
  .O(mux_o_3357),
  .I0(sdpb_inst_238_dout[26]),
  .I1(sdpb_inst_239_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3358 (
  .O(mux_o_3358),
  .I0(sdpb_inst_240_dout[26]),
  .I1(sdpb_inst_241_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3359 (
  .O(mux_o_3359),
  .I0(sdpb_inst_242_dout[26]),
  .I1(sdpb_inst_243_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3360 (
  .O(mux_o_3360),
  .I0(sdpb_inst_244_dout[26]),
  .I1(sdpb_inst_245_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3361 (
  .O(mux_o_3361),
  .I0(sdpb_inst_246_dout[26]),
  .I1(sdpb_inst_247_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3362 (
  .O(mux_o_3362),
  .I0(sdpb_inst_248_dout[26]),
  .I1(sdpb_inst_249_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3363 (
  .O(mux_o_3363),
  .I0(sdpb_inst_250_dout[26]),
  .I1(sdpb_inst_251_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3364 (
  .O(mux_o_3364),
  .I0(sdpb_inst_252_dout[26]),
  .I1(sdpb_inst_253_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3365 (
  .O(mux_o_3365),
  .I0(sdpb_inst_254_dout[26]),
  .I1(sdpb_inst_255_dout[26]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3366 (
  .O(mux_o_3366),
  .I0(mux_o_3302),
  .I1(mux_o_3303),
  .S0(dff_q_5)
);
MUX2 mux_inst_3367 (
  .O(mux_o_3367),
  .I0(mux_o_3304),
  .I1(mux_o_3305),
  .S0(dff_q_5)
);
MUX2 mux_inst_3368 (
  .O(mux_o_3368),
  .I0(mux_o_3306),
  .I1(mux_o_3307),
  .S0(dff_q_5)
);
MUX2 mux_inst_3369 (
  .O(mux_o_3369),
  .I0(mux_o_3308),
  .I1(mux_o_3309),
  .S0(dff_q_5)
);
MUX2 mux_inst_3370 (
  .O(mux_o_3370),
  .I0(mux_o_3310),
  .I1(mux_o_3311),
  .S0(dff_q_5)
);
MUX2 mux_inst_3371 (
  .O(mux_o_3371),
  .I0(mux_o_3312),
  .I1(mux_o_3313),
  .S0(dff_q_5)
);
MUX2 mux_inst_3372 (
  .O(mux_o_3372),
  .I0(mux_o_3314),
  .I1(mux_o_3315),
  .S0(dff_q_5)
);
MUX2 mux_inst_3373 (
  .O(mux_o_3373),
  .I0(mux_o_3316),
  .I1(mux_o_3317),
  .S0(dff_q_5)
);
MUX2 mux_inst_3374 (
  .O(mux_o_3374),
  .I0(mux_o_3318),
  .I1(mux_o_3319),
  .S0(dff_q_5)
);
MUX2 mux_inst_3375 (
  .O(mux_o_3375),
  .I0(mux_o_3320),
  .I1(mux_o_3321),
  .S0(dff_q_5)
);
MUX2 mux_inst_3376 (
  .O(mux_o_3376),
  .I0(mux_o_3322),
  .I1(mux_o_3323),
  .S0(dff_q_5)
);
MUX2 mux_inst_3377 (
  .O(mux_o_3377),
  .I0(mux_o_3324),
  .I1(mux_o_3325),
  .S0(dff_q_5)
);
MUX2 mux_inst_3378 (
  .O(mux_o_3378),
  .I0(mux_o_3326),
  .I1(mux_o_3327),
  .S0(dff_q_5)
);
MUX2 mux_inst_3379 (
  .O(mux_o_3379),
  .I0(mux_o_3328),
  .I1(mux_o_3329),
  .S0(dff_q_5)
);
MUX2 mux_inst_3380 (
  .O(mux_o_3380),
  .I0(mux_o_3330),
  .I1(mux_o_3331),
  .S0(dff_q_5)
);
MUX2 mux_inst_3381 (
  .O(mux_o_3381),
  .I0(mux_o_3332),
  .I1(mux_o_3333),
  .S0(dff_q_5)
);
MUX2 mux_inst_3382 (
  .O(mux_o_3382),
  .I0(mux_o_3334),
  .I1(mux_o_3335),
  .S0(dff_q_5)
);
MUX2 mux_inst_3383 (
  .O(mux_o_3383),
  .I0(mux_o_3336),
  .I1(mux_o_3337),
  .S0(dff_q_5)
);
MUX2 mux_inst_3384 (
  .O(mux_o_3384),
  .I0(mux_o_3338),
  .I1(mux_o_3339),
  .S0(dff_q_5)
);
MUX2 mux_inst_3385 (
  .O(mux_o_3385),
  .I0(mux_o_3340),
  .I1(mux_o_3341),
  .S0(dff_q_5)
);
MUX2 mux_inst_3386 (
  .O(mux_o_3386),
  .I0(mux_o_3342),
  .I1(mux_o_3343),
  .S0(dff_q_5)
);
MUX2 mux_inst_3387 (
  .O(mux_o_3387),
  .I0(mux_o_3344),
  .I1(mux_o_3345),
  .S0(dff_q_5)
);
MUX2 mux_inst_3388 (
  .O(mux_o_3388),
  .I0(mux_o_3346),
  .I1(mux_o_3347),
  .S0(dff_q_5)
);
MUX2 mux_inst_3389 (
  .O(mux_o_3389),
  .I0(mux_o_3348),
  .I1(mux_o_3349),
  .S0(dff_q_5)
);
MUX2 mux_inst_3390 (
  .O(mux_o_3390),
  .I0(mux_o_3350),
  .I1(mux_o_3351),
  .S0(dff_q_5)
);
MUX2 mux_inst_3391 (
  .O(mux_o_3391),
  .I0(mux_o_3352),
  .I1(mux_o_3353),
  .S0(dff_q_5)
);
MUX2 mux_inst_3392 (
  .O(mux_o_3392),
  .I0(mux_o_3354),
  .I1(mux_o_3355),
  .S0(dff_q_5)
);
MUX2 mux_inst_3393 (
  .O(mux_o_3393),
  .I0(mux_o_3356),
  .I1(mux_o_3357),
  .S0(dff_q_5)
);
MUX2 mux_inst_3394 (
  .O(mux_o_3394),
  .I0(mux_o_3358),
  .I1(mux_o_3359),
  .S0(dff_q_5)
);
MUX2 mux_inst_3395 (
  .O(mux_o_3395),
  .I0(mux_o_3360),
  .I1(mux_o_3361),
  .S0(dff_q_5)
);
MUX2 mux_inst_3396 (
  .O(mux_o_3396),
  .I0(mux_o_3362),
  .I1(mux_o_3363),
  .S0(dff_q_5)
);
MUX2 mux_inst_3397 (
  .O(mux_o_3397),
  .I0(mux_o_3364),
  .I1(mux_o_3365),
  .S0(dff_q_5)
);
MUX2 mux_inst_3398 (
  .O(mux_o_3398),
  .I0(mux_o_3366),
  .I1(mux_o_3367),
  .S0(dff_q_4)
);
MUX2 mux_inst_3399 (
  .O(mux_o_3399),
  .I0(mux_o_3368),
  .I1(mux_o_3369),
  .S0(dff_q_4)
);
MUX2 mux_inst_3400 (
  .O(mux_o_3400),
  .I0(mux_o_3370),
  .I1(mux_o_3371),
  .S0(dff_q_4)
);
MUX2 mux_inst_3401 (
  .O(mux_o_3401),
  .I0(mux_o_3372),
  .I1(mux_o_3373),
  .S0(dff_q_4)
);
MUX2 mux_inst_3402 (
  .O(mux_o_3402),
  .I0(mux_o_3374),
  .I1(mux_o_3375),
  .S0(dff_q_4)
);
MUX2 mux_inst_3403 (
  .O(mux_o_3403),
  .I0(mux_o_3376),
  .I1(mux_o_3377),
  .S0(dff_q_4)
);
MUX2 mux_inst_3404 (
  .O(mux_o_3404),
  .I0(mux_o_3378),
  .I1(mux_o_3379),
  .S0(dff_q_4)
);
MUX2 mux_inst_3405 (
  .O(mux_o_3405),
  .I0(mux_o_3380),
  .I1(mux_o_3381),
  .S0(dff_q_4)
);
MUX2 mux_inst_3406 (
  .O(mux_o_3406),
  .I0(mux_o_3382),
  .I1(mux_o_3383),
  .S0(dff_q_4)
);
MUX2 mux_inst_3407 (
  .O(mux_o_3407),
  .I0(mux_o_3384),
  .I1(mux_o_3385),
  .S0(dff_q_4)
);
MUX2 mux_inst_3408 (
  .O(mux_o_3408),
  .I0(mux_o_3386),
  .I1(mux_o_3387),
  .S0(dff_q_4)
);
MUX2 mux_inst_3409 (
  .O(mux_o_3409),
  .I0(mux_o_3388),
  .I1(mux_o_3389),
  .S0(dff_q_4)
);
MUX2 mux_inst_3410 (
  .O(mux_o_3410),
  .I0(mux_o_3390),
  .I1(mux_o_3391),
  .S0(dff_q_4)
);
MUX2 mux_inst_3411 (
  .O(mux_o_3411),
  .I0(mux_o_3392),
  .I1(mux_o_3393),
  .S0(dff_q_4)
);
MUX2 mux_inst_3412 (
  .O(mux_o_3412),
  .I0(mux_o_3394),
  .I1(mux_o_3395),
  .S0(dff_q_4)
);
MUX2 mux_inst_3413 (
  .O(mux_o_3413),
  .I0(mux_o_3396),
  .I1(mux_o_3397),
  .S0(dff_q_4)
);
MUX2 mux_inst_3414 (
  .O(mux_o_3414),
  .I0(mux_o_3398),
  .I1(mux_o_3399),
  .S0(dff_q_3)
);
MUX2 mux_inst_3415 (
  .O(mux_o_3415),
  .I0(mux_o_3400),
  .I1(mux_o_3401),
  .S0(dff_q_3)
);
MUX2 mux_inst_3416 (
  .O(mux_o_3416),
  .I0(mux_o_3402),
  .I1(mux_o_3403),
  .S0(dff_q_3)
);
MUX2 mux_inst_3417 (
  .O(mux_o_3417),
  .I0(mux_o_3404),
  .I1(mux_o_3405),
  .S0(dff_q_3)
);
MUX2 mux_inst_3418 (
  .O(mux_o_3418),
  .I0(mux_o_3406),
  .I1(mux_o_3407),
  .S0(dff_q_3)
);
MUX2 mux_inst_3419 (
  .O(mux_o_3419),
  .I0(mux_o_3408),
  .I1(mux_o_3409),
  .S0(dff_q_3)
);
MUX2 mux_inst_3420 (
  .O(mux_o_3420),
  .I0(mux_o_3410),
  .I1(mux_o_3411),
  .S0(dff_q_3)
);
MUX2 mux_inst_3421 (
  .O(mux_o_3421),
  .I0(mux_o_3412),
  .I1(mux_o_3413),
  .S0(dff_q_3)
);
MUX2 mux_inst_3422 (
  .O(mux_o_3422),
  .I0(mux_o_3414),
  .I1(mux_o_3415),
  .S0(dff_q_2)
);
MUX2 mux_inst_3423 (
  .O(mux_o_3423),
  .I0(mux_o_3416),
  .I1(mux_o_3417),
  .S0(dff_q_2)
);
MUX2 mux_inst_3424 (
  .O(mux_o_3424),
  .I0(mux_o_3418),
  .I1(mux_o_3419),
  .S0(dff_q_2)
);
MUX2 mux_inst_3425 (
  .O(mux_o_3425),
  .I0(mux_o_3420),
  .I1(mux_o_3421),
  .S0(dff_q_2)
);
MUX2 mux_inst_3426 (
  .O(mux_o_3426),
  .I0(mux_o_3422),
  .I1(mux_o_3423),
  .S0(dff_q_1)
);
MUX2 mux_inst_3427 (
  .O(mux_o_3427),
  .I0(mux_o_3424),
  .I1(mux_o_3425),
  .S0(dff_q_1)
);
MUX2 mux_inst_3428 (
  .O(dout[26]),
  .I0(mux_o_3426),
  .I1(mux_o_3427),
  .S0(dff_q_0)
);
MUX2 mux_inst_3429 (
  .O(mux_o_3429),
  .I0(sdpb_inst_128_dout[27]),
  .I1(sdpb_inst_129_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3430 (
  .O(mux_o_3430),
  .I0(sdpb_inst_130_dout[27]),
  .I1(sdpb_inst_131_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3431 (
  .O(mux_o_3431),
  .I0(sdpb_inst_132_dout[27]),
  .I1(sdpb_inst_133_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3432 (
  .O(mux_o_3432),
  .I0(sdpb_inst_134_dout[27]),
  .I1(sdpb_inst_135_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3433 (
  .O(mux_o_3433),
  .I0(sdpb_inst_136_dout[27]),
  .I1(sdpb_inst_137_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3434 (
  .O(mux_o_3434),
  .I0(sdpb_inst_138_dout[27]),
  .I1(sdpb_inst_139_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3435 (
  .O(mux_o_3435),
  .I0(sdpb_inst_140_dout[27]),
  .I1(sdpb_inst_141_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3436 (
  .O(mux_o_3436),
  .I0(sdpb_inst_142_dout[27]),
  .I1(sdpb_inst_143_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3437 (
  .O(mux_o_3437),
  .I0(sdpb_inst_144_dout[27]),
  .I1(sdpb_inst_145_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3438 (
  .O(mux_o_3438),
  .I0(sdpb_inst_146_dout[27]),
  .I1(sdpb_inst_147_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3439 (
  .O(mux_o_3439),
  .I0(sdpb_inst_148_dout[27]),
  .I1(sdpb_inst_149_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3440 (
  .O(mux_o_3440),
  .I0(sdpb_inst_150_dout[27]),
  .I1(sdpb_inst_151_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3441 (
  .O(mux_o_3441),
  .I0(sdpb_inst_152_dout[27]),
  .I1(sdpb_inst_153_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3442 (
  .O(mux_o_3442),
  .I0(sdpb_inst_154_dout[27]),
  .I1(sdpb_inst_155_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3443 (
  .O(mux_o_3443),
  .I0(sdpb_inst_156_dout[27]),
  .I1(sdpb_inst_157_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3444 (
  .O(mux_o_3444),
  .I0(sdpb_inst_158_dout[27]),
  .I1(sdpb_inst_159_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3445 (
  .O(mux_o_3445),
  .I0(sdpb_inst_160_dout[27]),
  .I1(sdpb_inst_161_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3446 (
  .O(mux_o_3446),
  .I0(sdpb_inst_162_dout[27]),
  .I1(sdpb_inst_163_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3447 (
  .O(mux_o_3447),
  .I0(sdpb_inst_164_dout[27]),
  .I1(sdpb_inst_165_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3448 (
  .O(mux_o_3448),
  .I0(sdpb_inst_166_dout[27]),
  .I1(sdpb_inst_167_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3449 (
  .O(mux_o_3449),
  .I0(sdpb_inst_168_dout[27]),
  .I1(sdpb_inst_169_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3450 (
  .O(mux_o_3450),
  .I0(sdpb_inst_170_dout[27]),
  .I1(sdpb_inst_171_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3451 (
  .O(mux_o_3451),
  .I0(sdpb_inst_172_dout[27]),
  .I1(sdpb_inst_173_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3452 (
  .O(mux_o_3452),
  .I0(sdpb_inst_174_dout[27]),
  .I1(sdpb_inst_175_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3453 (
  .O(mux_o_3453),
  .I0(sdpb_inst_176_dout[27]),
  .I1(sdpb_inst_177_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3454 (
  .O(mux_o_3454),
  .I0(sdpb_inst_178_dout[27]),
  .I1(sdpb_inst_179_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3455 (
  .O(mux_o_3455),
  .I0(sdpb_inst_180_dout[27]),
  .I1(sdpb_inst_181_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3456 (
  .O(mux_o_3456),
  .I0(sdpb_inst_182_dout[27]),
  .I1(sdpb_inst_183_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3457 (
  .O(mux_o_3457),
  .I0(sdpb_inst_184_dout[27]),
  .I1(sdpb_inst_185_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3458 (
  .O(mux_o_3458),
  .I0(sdpb_inst_186_dout[27]),
  .I1(sdpb_inst_187_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3459 (
  .O(mux_o_3459),
  .I0(sdpb_inst_188_dout[27]),
  .I1(sdpb_inst_189_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3460 (
  .O(mux_o_3460),
  .I0(sdpb_inst_190_dout[27]),
  .I1(sdpb_inst_191_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3461 (
  .O(mux_o_3461),
  .I0(sdpb_inst_192_dout[27]),
  .I1(sdpb_inst_193_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3462 (
  .O(mux_o_3462),
  .I0(sdpb_inst_194_dout[27]),
  .I1(sdpb_inst_195_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3463 (
  .O(mux_o_3463),
  .I0(sdpb_inst_196_dout[27]),
  .I1(sdpb_inst_197_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3464 (
  .O(mux_o_3464),
  .I0(sdpb_inst_198_dout[27]),
  .I1(sdpb_inst_199_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3465 (
  .O(mux_o_3465),
  .I0(sdpb_inst_200_dout[27]),
  .I1(sdpb_inst_201_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3466 (
  .O(mux_o_3466),
  .I0(sdpb_inst_202_dout[27]),
  .I1(sdpb_inst_203_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3467 (
  .O(mux_o_3467),
  .I0(sdpb_inst_204_dout[27]),
  .I1(sdpb_inst_205_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3468 (
  .O(mux_o_3468),
  .I0(sdpb_inst_206_dout[27]),
  .I1(sdpb_inst_207_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3469 (
  .O(mux_o_3469),
  .I0(sdpb_inst_208_dout[27]),
  .I1(sdpb_inst_209_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3470 (
  .O(mux_o_3470),
  .I0(sdpb_inst_210_dout[27]),
  .I1(sdpb_inst_211_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3471 (
  .O(mux_o_3471),
  .I0(sdpb_inst_212_dout[27]),
  .I1(sdpb_inst_213_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3472 (
  .O(mux_o_3472),
  .I0(sdpb_inst_214_dout[27]),
  .I1(sdpb_inst_215_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3473 (
  .O(mux_o_3473),
  .I0(sdpb_inst_216_dout[27]),
  .I1(sdpb_inst_217_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3474 (
  .O(mux_o_3474),
  .I0(sdpb_inst_218_dout[27]),
  .I1(sdpb_inst_219_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3475 (
  .O(mux_o_3475),
  .I0(sdpb_inst_220_dout[27]),
  .I1(sdpb_inst_221_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3476 (
  .O(mux_o_3476),
  .I0(sdpb_inst_222_dout[27]),
  .I1(sdpb_inst_223_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3477 (
  .O(mux_o_3477),
  .I0(sdpb_inst_224_dout[27]),
  .I1(sdpb_inst_225_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3478 (
  .O(mux_o_3478),
  .I0(sdpb_inst_226_dout[27]),
  .I1(sdpb_inst_227_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3479 (
  .O(mux_o_3479),
  .I0(sdpb_inst_228_dout[27]),
  .I1(sdpb_inst_229_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3480 (
  .O(mux_o_3480),
  .I0(sdpb_inst_230_dout[27]),
  .I1(sdpb_inst_231_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3481 (
  .O(mux_o_3481),
  .I0(sdpb_inst_232_dout[27]),
  .I1(sdpb_inst_233_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3482 (
  .O(mux_o_3482),
  .I0(sdpb_inst_234_dout[27]),
  .I1(sdpb_inst_235_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3483 (
  .O(mux_o_3483),
  .I0(sdpb_inst_236_dout[27]),
  .I1(sdpb_inst_237_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3484 (
  .O(mux_o_3484),
  .I0(sdpb_inst_238_dout[27]),
  .I1(sdpb_inst_239_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3485 (
  .O(mux_o_3485),
  .I0(sdpb_inst_240_dout[27]),
  .I1(sdpb_inst_241_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3486 (
  .O(mux_o_3486),
  .I0(sdpb_inst_242_dout[27]),
  .I1(sdpb_inst_243_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3487 (
  .O(mux_o_3487),
  .I0(sdpb_inst_244_dout[27]),
  .I1(sdpb_inst_245_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3488 (
  .O(mux_o_3488),
  .I0(sdpb_inst_246_dout[27]),
  .I1(sdpb_inst_247_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3489 (
  .O(mux_o_3489),
  .I0(sdpb_inst_248_dout[27]),
  .I1(sdpb_inst_249_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3490 (
  .O(mux_o_3490),
  .I0(sdpb_inst_250_dout[27]),
  .I1(sdpb_inst_251_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3491 (
  .O(mux_o_3491),
  .I0(sdpb_inst_252_dout[27]),
  .I1(sdpb_inst_253_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3492 (
  .O(mux_o_3492),
  .I0(sdpb_inst_254_dout[27]),
  .I1(sdpb_inst_255_dout[27]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3493 (
  .O(mux_o_3493),
  .I0(mux_o_3429),
  .I1(mux_o_3430),
  .S0(dff_q_5)
);
MUX2 mux_inst_3494 (
  .O(mux_o_3494),
  .I0(mux_o_3431),
  .I1(mux_o_3432),
  .S0(dff_q_5)
);
MUX2 mux_inst_3495 (
  .O(mux_o_3495),
  .I0(mux_o_3433),
  .I1(mux_o_3434),
  .S0(dff_q_5)
);
MUX2 mux_inst_3496 (
  .O(mux_o_3496),
  .I0(mux_o_3435),
  .I1(mux_o_3436),
  .S0(dff_q_5)
);
MUX2 mux_inst_3497 (
  .O(mux_o_3497),
  .I0(mux_o_3437),
  .I1(mux_o_3438),
  .S0(dff_q_5)
);
MUX2 mux_inst_3498 (
  .O(mux_o_3498),
  .I0(mux_o_3439),
  .I1(mux_o_3440),
  .S0(dff_q_5)
);
MUX2 mux_inst_3499 (
  .O(mux_o_3499),
  .I0(mux_o_3441),
  .I1(mux_o_3442),
  .S0(dff_q_5)
);
MUX2 mux_inst_3500 (
  .O(mux_o_3500),
  .I0(mux_o_3443),
  .I1(mux_o_3444),
  .S0(dff_q_5)
);
MUX2 mux_inst_3501 (
  .O(mux_o_3501),
  .I0(mux_o_3445),
  .I1(mux_o_3446),
  .S0(dff_q_5)
);
MUX2 mux_inst_3502 (
  .O(mux_o_3502),
  .I0(mux_o_3447),
  .I1(mux_o_3448),
  .S0(dff_q_5)
);
MUX2 mux_inst_3503 (
  .O(mux_o_3503),
  .I0(mux_o_3449),
  .I1(mux_o_3450),
  .S0(dff_q_5)
);
MUX2 mux_inst_3504 (
  .O(mux_o_3504),
  .I0(mux_o_3451),
  .I1(mux_o_3452),
  .S0(dff_q_5)
);
MUX2 mux_inst_3505 (
  .O(mux_o_3505),
  .I0(mux_o_3453),
  .I1(mux_o_3454),
  .S0(dff_q_5)
);
MUX2 mux_inst_3506 (
  .O(mux_o_3506),
  .I0(mux_o_3455),
  .I1(mux_o_3456),
  .S0(dff_q_5)
);
MUX2 mux_inst_3507 (
  .O(mux_o_3507),
  .I0(mux_o_3457),
  .I1(mux_o_3458),
  .S0(dff_q_5)
);
MUX2 mux_inst_3508 (
  .O(mux_o_3508),
  .I0(mux_o_3459),
  .I1(mux_o_3460),
  .S0(dff_q_5)
);
MUX2 mux_inst_3509 (
  .O(mux_o_3509),
  .I0(mux_o_3461),
  .I1(mux_o_3462),
  .S0(dff_q_5)
);
MUX2 mux_inst_3510 (
  .O(mux_o_3510),
  .I0(mux_o_3463),
  .I1(mux_o_3464),
  .S0(dff_q_5)
);
MUX2 mux_inst_3511 (
  .O(mux_o_3511),
  .I0(mux_o_3465),
  .I1(mux_o_3466),
  .S0(dff_q_5)
);
MUX2 mux_inst_3512 (
  .O(mux_o_3512),
  .I0(mux_o_3467),
  .I1(mux_o_3468),
  .S0(dff_q_5)
);
MUX2 mux_inst_3513 (
  .O(mux_o_3513),
  .I0(mux_o_3469),
  .I1(mux_o_3470),
  .S0(dff_q_5)
);
MUX2 mux_inst_3514 (
  .O(mux_o_3514),
  .I0(mux_o_3471),
  .I1(mux_o_3472),
  .S0(dff_q_5)
);
MUX2 mux_inst_3515 (
  .O(mux_o_3515),
  .I0(mux_o_3473),
  .I1(mux_o_3474),
  .S0(dff_q_5)
);
MUX2 mux_inst_3516 (
  .O(mux_o_3516),
  .I0(mux_o_3475),
  .I1(mux_o_3476),
  .S0(dff_q_5)
);
MUX2 mux_inst_3517 (
  .O(mux_o_3517),
  .I0(mux_o_3477),
  .I1(mux_o_3478),
  .S0(dff_q_5)
);
MUX2 mux_inst_3518 (
  .O(mux_o_3518),
  .I0(mux_o_3479),
  .I1(mux_o_3480),
  .S0(dff_q_5)
);
MUX2 mux_inst_3519 (
  .O(mux_o_3519),
  .I0(mux_o_3481),
  .I1(mux_o_3482),
  .S0(dff_q_5)
);
MUX2 mux_inst_3520 (
  .O(mux_o_3520),
  .I0(mux_o_3483),
  .I1(mux_o_3484),
  .S0(dff_q_5)
);
MUX2 mux_inst_3521 (
  .O(mux_o_3521),
  .I0(mux_o_3485),
  .I1(mux_o_3486),
  .S0(dff_q_5)
);
MUX2 mux_inst_3522 (
  .O(mux_o_3522),
  .I0(mux_o_3487),
  .I1(mux_o_3488),
  .S0(dff_q_5)
);
MUX2 mux_inst_3523 (
  .O(mux_o_3523),
  .I0(mux_o_3489),
  .I1(mux_o_3490),
  .S0(dff_q_5)
);
MUX2 mux_inst_3524 (
  .O(mux_o_3524),
  .I0(mux_o_3491),
  .I1(mux_o_3492),
  .S0(dff_q_5)
);
MUX2 mux_inst_3525 (
  .O(mux_o_3525),
  .I0(mux_o_3493),
  .I1(mux_o_3494),
  .S0(dff_q_4)
);
MUX2 mux_inst_3526 (
  .O(mux_o_3526),
  .I0(mux_o_3495),
  .I1(mux_o_3496),
  .S0(dff_q_4)
);
MUX2 mux_inst_3527 (
  .O(mux_o_3527),
  .I0(mux_o_3497),
  .I1(mux_o_3498),
  .S0(dff_q_4)
);
MUX2 mux_inst_3528 (
  .O(mux_o_3528),
  .I0(mux_o_3499),
  .I1(mux_o_3500),
  .S0(dff_q_4)
);
MUX2 mux_inst_3529 (
  .O(mux_o_3529),
  .I0(mux_o_3501),
  .I1(mux_o_3502),
  .S0(dff_q_4)
);
MUX2 mux_inst_3530 (
  .O(mux_o_3530),
  .I0(mux_o_3503),
  .I1(mux_o_3504),
  .S0(dff_q_4)
);
MUX2 mux_inst_3531 (
  .O(mux_o_3531),
  .I0(mux_o_3505),
  .I1(mux_o_3506),
  .S0(dff_q_4)
);
MUX2 mux_inst_3532 (
  .O(mux_o_3532),
  .I0(mux_o_3507),
  .I1(mux_o_3508),
  .S0(dff_q_4)
);
MUX2 mux_inst_3533 (
  .O(mux_o_3533),
  .I0(mux_o_3509),
  .I1(mux_o_3510),
  .S0(dff_q_4)
);
MUX2 mux_inst_3534 (
  .O(mux_o_3534),
  .I0(mux_o_3511),
  .I1(mux_o_3512),
  .S0(dff_q_4)
);
MUX2 mux_inst_3535 (
  .O(mux_o_3535),
  .I0(mux_o_3513),
  .I1(mux_o_3514),
  .S0(dff_q_4)
);
MUX2 mux_inst_3536 (
  .O(mux_o_3536),
  .I0(mux_o_3515),
  .I1(mux_o_3516),
  .S0(dff_q_4)
);
MUX2 mux_inst_3537 (
  .O(mux_o_3537),
  .I0(mux_o_3517),
  .I1(mux_o_3518),
  .S0(dff_q_4)
);
MUX2 mux_inst_3538 (
  .O(mux_o_3538),
  .I0(mux_o_3519),
  .I1(mux_o_3520),
  .S0(dff_q_4)
);
MUX2 mux_inst_3539 (
  .O(mux_o_3539),
  .I0(mux_o_3521),
  .I1(mux_o_3522),
  .S0(dff_q_4)
);
MUX2 mux_inst_3540 (
  .O(mux_o_3540),
  .I0(mux_o_3523),
  .I1(mux_o_3524),
  .S0(dff_q_4)
);
MUX2 mux_inst_3541 (
  .O(mux_o_3541),
  .I0(mux_o_3525),
  .I1(mux_o_3526),
  .S0(dff_q_3)
);
MUX2 mux_inst_3542 (
  .O(mux_o_3542),
  .I0(mux_o_3527),
  .I1(mux_o_3528),
  .S0(dff_q_3)
);
MUX2 mux_inst_3543 (
  .O(mux_o_3543),
  .I0(mux_o_3529),
  .I1(mux_o_3530),
  .S0(dff_q_3)
);
MUX2 mux_inst_3544 (
  .O(mux_o_3544),
  .I0(mux_o_3531),
  .I1(mux_o_3532),
  .S0(dff_q_3)
);
MUX2 mux_inst_3545 (
  .O(mux_o_3545),
  .I0(mux_o_3533),
  .I1(mux_o_3534),
  .S0(dff_q_3)
);
MUX2 mux_inst_3546 (
  .O(mux_o_3546),
  .I0(mux_o_3535),
  .I1(mux_o_3536),
  .S0(dff_q_3)
);
MUX2 mux_inst_3547 (
  .O(mux_o_3547),
  .I0(mux_o_3537),
  .I1(mux_o_3538),
  .S0(dff_q_3)
);
MUX2 mux_inst_3548 (
  .O(mux_o_3548),
  .I0(mux_o_3539),
  .I1(mux_o_3540),
  .S0(dff_q_3)
);
MUX2 mux_inst_3549 (
  .O(mux_o_3549),
  .I0(mux_o_3541),
  .I1(mux_o_3542),
  .S0(dff_q_2)
);
MUX2 mux_inst_3550 (
  .O(mux_o_3550),
  .I0(mux_o_3543),
  .I1(mux_o_3544),
  .S0(dff_q_2)
);
MUX2 mux_inst_3551 (
  .O(mux_o_3551),
  .I0(mux_o_3545),
  .I1(mux_o_3546),
  .S0(dff_q_2)
);
MUX2 mux_inst_3552 (
  .O(mux_o_3552),
  .I0(mux_o_3547),
  .I1(mux_o_3548),
  .S0(dff_q_2)
);
MUX2 mux_inst_3553 (
  .O(mux_o_3553),
  .I0(mux_o_3549),
  .I1(mux_o_3550),
  .S0(dff_q_1)
);
MUX2 mux_inst_3554 (
  .O(mux_o_3554),
  .I0(mux_o_3551),
  .I1(mux_o_3552),
  .S0(dff_q_1)
);
MUX2 mux_inst_3555 (
  .O(dout[27]),
  .I0(mux_o_3553),
  .I1(mux_o_3554),
  .S0(dff_q_0)
);
MUX2 mux_inst_3556 (
  .O(mux_o_3556),
  .I0(sdpb_inst_128_dout[28]),
  .I1(sdpb_inst_129_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3557 (
  .O(mux_o_3557),
  .I0(sdpb_inst_130_dout[28]),
  .I1(sdpb_inst_131_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3558 (
  .O(mux_o_3558),
  .I0(sdpb_inst_132_dout[28]),
  .I1(sdpb_inst_133_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3559 (
  .O(mux_o_3559),
  .I0(sdpb_inst_134_dout[28]),
  .I1(sdpb_inst_135_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3560 (
  .O(mux_o_3560),
  .I0(sdpb_inst_136_dout[28]),
  .I1(sdpb_inst_137_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3561 (
  .O(mux_o_3561),
  .I0(sdpb_inst_138_dout[28]),
  .I1(sdpb_inst_139_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3562 (
  .O(mux_o_3562),
  .I0(sdpb_inst_140_dout[28]),
  .I1(sdpb_inst_141_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3563 (
  .O(mux_o_3563),
  .I0(sdpb_inst_142_dout[28]),
  .I1(sdpb_inst_143_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3564 (
  .O(mux_o_3564),
  .I0(sdpb_inst_144_dout[28]),
  .I1(sdpb_inst_145_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3565 (
  .O(mux_o_3565),
  .I0(sdpb_inst_146_dout[28]),
  .I1(sdpb_inst_147_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3566 (
  .O(mux_o_3566),
  .I0(sdpb_inst_148_dout[28]),
  .I1(sdpb_inst_149_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3567 (
  .O(mux_o_3567),
  .I0(sdpb_inst_150_dout[28]),
  .I1(sdpb_inst_151_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3568 (
  .O(mux_o_3568),
  .I0(sdpb_inst_152_dout[28]),
  .I1(sdpb_inst_153_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3569 (
  .O(mux_o_3569),
  .I0(sdpb_inst_154_dout[28]),
  .I1(sdpb_inst_155_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3570 (
  .O(mux_o_3570),
  .I0(sdpb_inst_156_dout[28]),
  .I1(sdpb_inst_157_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3571 (
  .O(mux_o_3571),
  .I0(sdpb_inst_158_dout[28]),
  .I1(sdpb_inst_159_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3572 (
  .O(mux_o_3572),
  .I0(sdpb_inst_160_dout[28]),
  .I1(sdpb_inst_161_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3573 (
  .O(mux_o_3573),
  .I0(sdpb_inst_162_dout[28]),
  .I1(sdpb_inst_163_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3574 (
  .O(mux_o_3574),
  .I0(sdpb_inst_164_dout[28]),
  .I1(sdpb_inst_165_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3575 (
  .O(mux_o_3575),
  .I0(sdpb_inst_166_dout[28]),
  .I1(sdpb_inst_167_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3576 (
  .O(mux_o_3576),
  .I0(sdpb_inst_168_dout[28]),
  .I1(sdpb_inst_169_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3577 (
  .O(mux_o_3577),
  .I0(sdpb_inst_170_dout[28]),
  .I1(sdpb_inst_171_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3578 (
  .O(mux_o_3578),
  .I0(sdpb_inst_172_dout[28]),
  .I1(sdpb_inst_173_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3579 (
  .O(mux_o_3579),
  .I0(sdpb_inst_174_dout[28]),
  .I1(sdpb_inst_175_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3580 (
  .O(mux_o_3580),
  .I0(sdpb_inst_176_dout[28]),
  .I1(sdpb_inst_177_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3581 (
  .O(mux_o_3581),
  .I0(sdpb_inst_178_dout[28]),
  .I1(sdpb_inst_179_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3582 (
  .O(mux_o_3582),
  .I0(sdpb_inst_180_dout[28]),
  .I1(sdpb_inst_181_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3583 (
  .O(mux_o_3583),
  .I0(sdpb_inst_182_dout[28]),
  .I1(sdpb_inst_183_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3584 (
  .O(mux_o_3584),
  .I0(sdpb_inst_184_dout[28]),
  .I1(sdpb_inst_185_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3585 (
  .O(mux_o_3585),
  .I0(sdpb_inst_186_dout[28]),
  .I1(sdpb_inst_187_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3586 (
  .O(mux_o_3586),
  .I0(sdpb_inst_188_dout[28]),
  .I1(sdpb_inst_189_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3587 (
  .O(mux_o_3587),
  .I0(sdpb_inst_190_dout[28]),
  .I1(sdpb_inst_191_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3588 (
  .O(mux_o_3588),
  .I0(sdpb_inst_192_dout[28]),
  .I1(sdpb_inst_193_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3589 (
  .O(mux_o_3589),
  .I0(sdpb_inst_194_dout[28]),
  .I1(sdpb_inst_195_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3590 (
  .O(mux_o_3590),
  .I0(sdpb_inst_196_dout[28]),
  .I1(sdpb_inst_197_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3591 (
  .O(mux_o_3591),
  .I0(sdpb_inst_198_dout[28]),
  .I1(sdpb_inst_199_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3592 (
  .O(mux_o_3592),
  .I0(sdpb_inst_200_dout[28]),
  .I1(sdpb_inst_201_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3593 (
  .O(mux_o_3593),
  .I0(sdpb_inst_202_dout[28]),
  .I1(sdpb_inst_203_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3594 (
  .O(mux_o_3594),
  .I0(sdpb_inst_204_dout[28]),
  .I1(sdpb_inst_205_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3595 (
  .O(mux_o_3595),
  .I0(sdpb_inst_206_dout[28]),
  .I1(sdpb_inst_207_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3596 (
  .O(mux_o_3596),
  .I0(sdpb_inst_208_dout[28]),
  .I1(sdpb_inst_209_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3597 (
  .O(mux_o_3597),
  .I0(sdpb_inst_210_dout[28]),
  .I1(sdpb_inst_211_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3598 (
  .O(mux_o_3598),
  .I0(sdpb_inst_212_dout[28]),
  .I1(sdpb_inst_213_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3599 (
  .O(mux_o_3599),
  .I0(sdpb_inst_214_dout[28]),
  .I1(sdpb_inst_215_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3600 (
  .O(mux_o_3600),
  .I0(sdpb_inst_216_dout[28]),
  .I1(sdpb_inst_217_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3601 (
  .O(mux_o_3601),
  .I0(sdpb_inst_218_dout[28]),
  .I1(sdpb_inst_219_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3602 (
  .O(mux_o_3602),
  .I0(sdpb_inst_220_dout[28]),
  .I1(sdpb_inst_221_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3603 (
  .O(mux_o_3603),
  .I0(sdpb_inst_222_dout[28]),
  .I1(sdpb_inst_223_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3604 (
  .O(mux_o_3604),
  .I0(sdpb_inst_224_dout[28]),
  .I1(sdpb_inst_225_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3605 (
  .O(mux_o_3605),
  .I0(sdpb_inst_226_dout[28]),
  .I1(sdpb_inst_227_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3606 (
  .O(mux_o_3606),
  .I0(sdpb_inst_228_dout[28]),
  .I1(sdpb_inst_229_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3607 (
  .O(mux_o_3607),
  .I0(sdpb_inst_230_dout[28]),
  .I1(sdpb_inst_231_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3608 (
  .O(mux_o_3608),
  .I0(sdpb_inst_232_dout[28]),
  .I1(sdpb_inst_233_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3609 (
  .O(mux_o_3609),
  .I0(sdpb_inst_234_dout[28]),
  .I1(sdpb_inst_235_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3610 (
  .O(mux_o_3610),
  .I0(sdpb_inst_236_dout[28]),
  .I1(sdpb_inst_237_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3611 (
  .O(mux_o_3611),
  .I0(sdpb_inst_238_dout[28]),
  .I1(sdpb_inst_239_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3612 (
  .O(mux_o_3612),
  .I0(sdpb_inst_240_dout[28]),
  .I1(sdpb_inst_241_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3613 (
  .O(mux_o_3613),
  .I0(sdpb_inst_242_dout[28]),
  .I1(sdpb_inst_243_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3614 (
  .O(mux_o_3614),
  .I0(sdpb_inst_244_dout[28]),
  .I1(sdpb_inst_245_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3615 (
  .O(mux_o_3615),
  .I0(sdpb_inst_246_dout[28]),
  .I1(sdpb_inst_247_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3616 (
  .O(mux_o_3616),
  .I0(sdpb_inst_248_dout[28]),
  .I1(sdpb_inst_249_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3617 (
  .O(mux_o_3617),
  .I0(sdpb_inst_250_dout[28]),
  .I1(sdpb_inst_251_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3618 (
  .O(mux_o_3618),
  .I0(sdpb_inst_252_dout[28]),
  .I1(sdpb_inst_253_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3619 (
  .O(mux_o_3619),
  .I0(sdpb_inst_254_dout[28]),
  .I1(sdpb_inst_255_dout[28]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3620 (
  .O(mux_o_3620),
  .I0(mux_o_3556),
  .I1(mux_o_3557),
  .S0(dff_q_5)
);
MUX2 mux_inst_3621 (
  .O(mux_o_3621),
  .I0(mux_o_3558),
  .I1(mux_o_3559),
  .S0(dff_q_5)
);
MUX2 mux_inst_3622 (
  .O(mux_o_3622),
  .I0(mux_o_3560),
  .I1(mux_o_3561),
  .S0(dff_q_5)
);
MUX2 mux_inst_3623 (
  .O(mux_o_3623),
  .I0(mux_o_3562),
  .I1(mux_o_3563),
  .S0(dff_q_5)
);
MUX2 mux_inst_3624 (
  .O(mux_o_3624),
  .I0(mux_o_3564),
  .I1(mux_o_3565),
  .S0(dff_q_5)
);
MUX2 mux_inst_3625 (
  .O(mux_o_3625),
  .I0(mux_o_3566),
  .I1(mux_o_3567),
  .S0(dff_q_5)
);
MUX2 mux_inst_3626 (
  .O(mux_o_3626),
  .I0(mux_o_3568),
  .I1(mux_o_3569),
  .S0(dff_q_5)
);
MUX2 mux_inst_3627 (
  .O(mux_o_3627),
  .I0(mux_o_3570),
  .I1(mux_o_3571),
  .S0(dff_q_5)
);
MUX2 mux_inst_3628 (
  .O(mux_o_3628),
  .I0(mux_o_3572),
  .I1(mux_o_3573),
  .S0(dff_q_5)
);
MUX2 mux_inst_3629 (
  .O(mux_o_3629),
  .I0(mux_o_3574),
  .I1(mux_o_3575),
  .S0(dff_q_5)
);
MUX2 mux_inst_3630 (
  .O(mux_o_3630),
  .I0(mux_o_3576),
  .I1(mux_o_3577),
  .S0(dff_q_5)
);
MUX2 mux_inst_3631 (
  .O(mux_o_3631),
  .I0(mux_o_3578),
  .I1(mux_o_3579),
  .S0(dff_q_5)
);
MUX2 mux_inst_3632 (
  .O(mux_o_3632),
  .I0(mux_o_3580),
  .I1(mux_o_3581),
  .S0(dff_q_5)
);
MUX2 mux_inst_3633 (
  .O(mux_o_3633),
  .I0(mux_o_3582),
  .I1(mux_o_3583),
  .S0(dff_q_5)
);
MUX2 mux_inst_3634 (
  .O(mux_o_3634),
  .I0(mux_o_3584),
  .I1(mux_o_3585),
  .S0(dff_q_5)
);
MUX2 mux_inst_3635 (
  .O(mux_o_3635),
  .I0(mux_o_3586),
  .I1(mux_o_3587),
  .S0(dff_q_5)
);
MUX2 mux_inst_3636 (
  .O(mux_o_3636),
  .I0(mux_o_3588),
  .I1(mux_o_3589),
  .S0(dff_q_5)
);
MUX2 mux_inst_3637 (
  .O(mux_o_3637),
  .I0(mux_o_3590),
  .I1(mux_o_3591),
  .S0(dff_q_5)
);
MUX2 mux_inst_3638 (
  .O(mux_o_3638),
  .I0(mux_o_3592),
  .I1(mux_o_3593),
  .S0(dff_q_5)
);
MUX2 mux_inst_3639 (
  .O(mux_o_3639),
  .I0(mux_o_3594),
  .I1(mux_o_3595),
  .S0(dff_q_5)
);
MUX2 mux_inst_3640 (
  .O(mux_o_3640),
  .I0(mux_o_3596),
  .I1(mux_o_3597),
  .S0(dff_q_5)
);
MUX2 mux_inst_3641 (
  .O(mux_o_3641),
  .I0(mux_o_3598),
  .I1(mux_o_3599),
  .S0(dff_q_5)
);
MUX2 mux_inst_3642 (
  .O(mux_o_3642),
  .I0(mux_o_3600),
  .I1(mux_o_3601),
  .S0(dff_q_5)
);
MUX2 mux_inst_3643 (
  .O(mux_o_3643),
  .I0(mux_o_3602),
  .I1(mux_o_3603),
  .S0(dff_q_5)
);
MUX2 mux_inst_3644 (
  .O(mux_o_3644),
  .I0(mux_o_3604),
  .I1(mux_o_3605),
  .S0(dff_q_5)
);
MUX2 mux_inst_3645 (
  .O(mux_o_3645),
  .I0(mux_o_3606),
  .I1(mux_o_3607),
  .S0(dff_q_5)
);
MUX2 mux_inst_3646 (
  .O(mux_o_3646),
  .I0(mux_o_3608),
  .I1(mux_o_3609),
  .S0(dff_q_5)
);
MUX2 mux_inst_3647 (
  .O(mux_o_3647),
  .I0(mux_o_3610),
  .I1(mux_o_3611),
  .S0(dff_q_5)
);
MUX2 mux_inst_3648 (
  .O(mux_o_3648),
  .I0(mux_o_3612),
  .I1(mux_o_3613),
  .S0(dff_q_5)
);
MUX2 mux_inst_3649 (
  .O(mux_o_3649),
  .I0(mux_o_3614),
  .I1(mux_o_3615),
  .S0(dff_q_5)
);
MUX2 mux_inst_3650 (
  .O(mux_o_3650),
  .I0(mux_o_3616),
  .I1(mux_o_3617),
  .S0(dff_q_5)
);
MUX2 mux_inst_3651 (
  .O(mux_o_3651),
  .I0(mux_o_3618),
  .I1(mux_o_3619),
  .S0(dff_q_5)
);
MUX2 mux_inst_3652 (
  .O(mux_o_3652),
  .I0(mux_o_3620),
  .I1(mux_o_3621),
  .S0(dff_q_4)
);
MUX2 mux_inst_3653 (
  .O(mux_o_3653),
  .I0(mux_o_3622),
  .I1(mux_o_3623),
  .S0(dff_q_4)
);
MUX2 mux_inst_3654 (
  .O(mux_o_3654),
  .I0(mux_o_3624),
  .I1(mux_o_3625),
  .S0(dff_q_4)
);
MUX2 mux_inst_3655 (
  .O(mux_o_3655),
  .I0(mux_o_3626),
  .I1(mux_o_3627),
  .S0(dff_q_4)
);
MUX2 mux_inst_3656 (
  .O(mux_o_3656),
  .I0(mux_o_3628),
  .I1(mux_o_3629),
  .S0(dff_q_4)
);
MUX2 mux_inst_3657 (
  .O(mux_o_3657),
  .I0(mux_o_3630),
  .I1(mux_o_3631),
  .S0(dff_q_4)
);
MUX2 mux_inst_3658 (
  .O(mux_o_3658),
  .I0(mux_o_3632),
  .I1(mux_o_3633),
  .S0(dff_q_4)
);
MUX2 mux_inst_3659 (
  .O(mux_o_3659),
  .I0(mux_o_3634),
  .I1(mux_o_3635),
  .S0(dff_q_4)
);
MUX2 mux_inst_3660 (
  .O(mux_o_3660),
  .I0(mux_o_3636),
  .I1(mux_o_3637),
  .S0(dff_q_4)
);
MUX2 mux_inst_3661 (
  .O(mux_o_3661),
  .I0(mux_o_3638),
  .I1(mux_o_3639),
  .S0(dff_q_4)
);
MUX2 mux_inst_3662 (
  .O(mux_o_3662),
  .I0(mux_o_3640),
  .I1(mux_o_3641),
  .S0(dff_q_4)
);
MUX2 mux_inst_3663 (
  .O(mux_o_3663),
  .I0(mux_o_3642),
  .I1(mux_o_3643),
  .S0(dff_q_4)
);
MUX2 mux_inst_3664 (
  .O(mux_o_3664),
  .I0(mux_o_3644),
  .I1(mux_o_3645),
  .S0(dff_q_4)
);
MUX2 mux_inst_3665 (
  .O(mux_o_3665),
  .I0(mux_o_3646),
  .I1(mux_o_3647),
  .S0(dff_q_4)
);
MUX2 mux_inst_3666 (
  .O(mux_o_3666),
  .I0(mux_o_3648),
  .I1(mux_o_3649),
  .S0(dff_q_4)
);
MUX2 mux_inst_3667 (
  .O(mux_o_3667),
  .I0(mux_o_3650),
  .I1(mux_o_3651),
  .S0(dff_q_4)
);
MUX2 mux_inst_3668 (
  .O(mux_o_3668),
  .I0(mux_o_3652),
  .I1(mux_o_3653),
  .S0(dff_q_3)
);
MUX2 mux_inst_3669 (
  .O(mux_o_3669),
  .I0(mux_o_3654),
  .I1(mux_o_3655),
  .S0(dff_q_3)
);
MUX2 mux_inst_3670 (
  .O(mux_o_3670),
  .I0(mux_o_3656),
  .I1(mux_o_3657),
  .S0(dff_q_3)
);
MUX2 mux_inst_3671 (
  .O(mux_o_3671),
  .I0(mux_o_3658),
  .I1(mux_o_3659),
  .S0(dff_q_3)
);
MUX2 mux_inst_3672 (
  .O(mux_o_3672),
  .I0(mux_o_3660),
  .I1(mux_o_3661),
  .S0(dff_q_3)
);
MUX2 mux_inst_3673 (
  .O(mux_o_3673),
  .I0(mux_o_3662),
  .I1(mux_o_3663),
  .S0(dff_q_3)
);
MUX2 mux_inst_3674 (
  .O(mux_o_3674),
  .I0(mux_o_3664),
  .I1(mux_o_3665),
  .S0(dff_q_3)
);
MUX2 mux_inst_3675 (
  .O(mux_o_3675),
  .I0(mux_o_3666),
  .I1(mux_o_3667),
  .S0(dff_q_3)
);
MUX2 mux_inst_3676 (
  .O(mux_o_3676),
  .I0(mux_o_3668),
  .I1(mux_o_3669),
  .S0(dff_q_2)
);
MUX2 mux_inst_3677 (
  .O(mux_o_3677),
  .I0(mux_o_3670),
  .I1(mux_o_3671),
  .S0(dff_q_2)
);
MUX2 mux_inst_3678 (
  .O(mux_o_3678),
  .I0(mux_o_3672),
  .I1(mux_o_3673),
  .S0(dff_q_2)
);
MUX2 mux_inst_3679 (
  .O(mux_o_3679),
  .I0(mux_o_3674),
  .I1(mux_o_3675),
  .S0(dff_q_2)
);
MUX2 mux_inst_3680 (
  .O(mux_o_3680),
  .I0(mux_o_3676),
  .I1(mux_o_3677),
  .S0(dff_q_1)
);
MUX2 mux_inst_3681 (
  .O(mux_o_3681),
  .I0(mux_o_3678),
  .I1(mux_o_3679),
  .S0(dff_q_1)
);
MUX2 mux_inst_3682 (
  .O(dout[28]),
  .I0(mux_o_3680),
  .I1(mux_o_3681),
  .S0(dff_q_0)
);
MUX2 mux_inst_3683 (
  .O(mux_o_3683),
  .I0(sdpb_inst_128_dout[29]),
  .I1(sdpb_inst_129_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3684 (
  .O(mux_o_3684),
  .I0(sdpb_inst_130_dout[29]),
  .I1(sdpb_inst_131_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3685 (
  .O(mux_o_3685),
  .I0(sdpb_inst_132_dout[29]),
  .I1(sdpb_inst_133_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3686 (
  .O(mux_o_3686),
  .I0(sdpb_inst_134_dout[29]),
  .I1(sdpb_inst_135_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3687 (
  .O(mux_o_3687),
  .I0(sdpb_inst_136_dout[29]),
  .I1(sdpb_inst_137_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3688 (
  .O(mux_o_3688),
  .I0(sdpb_inst_138_dout[29]),
  .I1(sdpb_inst_139_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3689 (
  .O(mux_o_3689),
  .I0(sdpb_inst_140_dout[29]),
  .I1(sdpb_inst_141_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3690 (
  .O(mux_o_3690),
  .I0(sdpb_inst_142_dout[29]),
  .I1(sdpb_inst_143_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3691 (
  .O(mux_o_3691),
  .I0(sdpb_inst_144_dout[29]),
  .I1(sdpb_inst_145_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3692 (
  .O(mux_o_3692),
  .I0(sdpb_inst_146_dout[29]),
  .I1(sdpb_inst_147_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3693 (
  .O(mux_o_3693),
  .I0(sdpb_inst_148_dout[29]),
  .I1(sdpb_inst_149_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3694 (
  .O(mux_o_3694),
  .I0(sdpb_inst_150_dout[29]),
  .I1(sdpb_inst_151_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3695 (
  .O(mux_o_3695),
  .I0(sdpb_inst_152_dout[29]),
  .I1(sdpb_inst_153_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3696 (
  .O(mux_o_3696),
  .I0(sdpb_inst_154_dout[29]),
  .I1(sdpb_inst_155_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3697 (
  .O(mux_o_3697),
  .I0(sdpb_inst_156_dout[29]),
  .I1(sdpb_inst_157_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3698 (
  .O(mux_o_3698),
  .I0(sdpb_inst_158_dout[29]),
  .I1(sdpb_inst_159_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3699 (
  .O(mux_o_3699),
  .I0(sdpb_inst_160_dout[29]),
  .I1(sdpb_inst_161_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3700 (
  .O(mux_o_3700),
  .I0(sdpb_inst_162_dout[29]),
  .I1(sdpb_inst_163_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3701 (
  .O(mux_o_3701),
  .I0(sdpb_inst_164_dout[29]),
  .I1(sdpb_inst_165_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3702 (
  .O(mux_o_3702),
  .I0(sdpb_inst_166_dout[29]),
  .I1(sdpb_inst_167_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3703 (
  .O(mux_o_3703),
  .I0(sdpb_inst_168_dout[29]),
  .I1(sdpb_inst_169_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3704 (
  .O(mux_o_3704),
  .I0(sdpb_inst_170_dout[29]),
  .I1(sdpb_inst_171_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3705 (
  .O(mux_o_3705),
  .I0(sdpb_inst_172_dout[29]),
  .I1(sdpb_inst_173_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3706 (
  .O(mux_o_3706),
  .I0(sdpb_inst_174_dout[29]),
  .I1(sdpb_inst_175_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3707 (
  .O(mux_o_3707),
  .I0(sdpb_inst_176_dout[29]),
  .I1(sdpb_inst_177_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3708 (
  .O(mux_o_3708),
  .I0(sdpb_inst_178_dout[29]),
  .I1(sdpb_inst_179_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3709 (
  .O(mux_o_3709),
  .I0(sdpb_inst_180_dout[29]),
  .I1(sdpb_inst_181_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3710 (
  .O(mux_o_3710),
  .I0(sdpb_inst_182_dout[29]),
  .I1(sdpb_inst_183_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3711 (
  .O(mux_o_3711),
  .I0(sdpb_inst_184_dout[29]),
  .I1(sdpb_inst_185_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3712 (
  .O(mux_o_3712),
  .I0(sdpb_inst_186_dout[29]),
  .I1(sdpb_inst_187_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3713 (
  .O(mux_o_3713),
  .I0(sdpb_inst_188_dout[29]),
  .I1(sdpb_inst_189_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3714 (
  .O(mux_o_3714),
  .I0(sdpb_inst_190_dout[29]),
  .I1(sdpb_inst_191_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3715 (
  .O(mux_o_3715),
  .I0(sdpb_inst_192_dout[29]),
  .I1(sdpb_inst_193_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3716 (
  .O(mux_o_3716),
  .I0(sdpb_inst_194_dout[29]),
  .I1(sdpb_inst_195_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3717 (
  .O(mux_o_3717),
  .I0(sdpb_inst_196_dout[29]),
  .I1(sdpb_inst_197_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3718 (
  .O(mux_o_3718),
  .I0(sdpb_inst_198_dout[29]),
  .I1(sdpb_inst_199_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3719 (
  .O(mux_o_3719),
  .I0(sdpb_inst_200_dout[29]),
  .I1(sdpb_inst_201_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3720 (
  .O(mux_o_3720),
  .I0(sdpb_inst_202_dout[29]),
  .I1(sdpb_inst_203_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3721 (
  .O(mux_o_3721),
  .I0(sdpb_inst_204_dout[29]),
  .I1(sdpb_inst_205_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3722 (
  .O(mux_o_3722),
  .I0(sdpb_inst_206_dout[29]),
  .I1(sdpb_inst_207_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3723 (
  .O(mux_o_3723),
  .I0(sdpb_inst_208_dout[29]),
  .I1(sdpb_inst_209_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3724 (
  .O(mux_o_3724),
  .I0(sdpb_inst_210_dout[29]),
  .I1(sdpb_inst_211_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3725 (
  .O(mux_o_3725),
  .I0(sdpb_inst_212_dout[29]),
  .I1(sdpb_inst_213_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3726 (
  .O(mux_o_3726),
  .I0(sdpb_inst_214_dout[29]),
  .I1(sdpb_inst_215_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3727 (
  .O(mux_o_3727),
  .I0(sdpb_inst_216_dout[29]),
  .I1(sdpb_inst_217_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3728 (
  .O(mux_o_3728),
  .I0(sdpb_inst_218_dout[29]),
  .I1(sdpb_inst_219_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3729 (
  .O(mux_o_3729),
  .I0(sdpb_inst_220_dout[29]),
  .I1(sdpb_inst_221_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3730 (
  .O(mux_o_3730),
  .I0(sdpb_inst_222_dout[29]),
  .I1(sdpb_inst_223_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3731 (
  .O(mux_o_3731),
  .I0(sdpb_inst_224_dout[29]),
  .I1(sdpb_inst_225_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3732 (
  .O(mux_o_3732),
  .I0(sdpb_inst_226_dout[29]),
  .I1(sdpb_inst_227_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3733 (
  .O(mux_o_3733),
  .I0(sdpb_inst_228_dout[29]),
  .I1(sdpb_inst_229_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3734 (
  .O(mux_o_3734),
  .I0(sdpb_inst_230_dout[29]),
  .I1(sdpb_inst_231_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3735 (
  .O(mux_o_3735),
  .I0(sdpb_inst_232_dout[29]),
  .I1(sdpb_inst_233_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3736 (
  .O(mux_o_3736),
  .I0(sdpb_inst_234_dout[29]),
  .I1(sdpb_inst_235_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3737 (
  .O(mux_o_3737),
  .I0(sdpb_inst_236_dout[29]),
  .I1(sdpb_inst_237_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3738 (
  .O(mux_o_3738),
  .I0(sdpb_inst_238_dout[29]),
  .I1(sdpb_inst_239_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3739 (
  .O(mux_o_3739),
  .I0(sdpb_inst_240_dout[29]),
  .I1(sdpb_inst_241_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3740 (
  .O(mux_o_3740),
  .I0(sdpb_inst_242_dout[29]),
  .I1(sdpb_inst_243_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3741 (
  .O(mux_o_3741),
  .I0(sdpb_inst_244_dout[29]),
  .I1(sdpb_inst_245_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3742 (
  .O(mux_o_3742),
  .I0(sdpb_inst_246_dout[29]),
  .I1(sdpb_inst_247_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3743 (
  .O(mux_o_3743),
  .I0(sdpb_inst_248_dout[29]),
  .I1(sdpb_inst_249_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3744 (
  .O(mux_o_3744),
  .I0(sdpb_inst_250_dout[29]),
  .I1(sdpb_inst_251_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3745 (
  .O(mux_o_3745),
  .I0(sdpb_inst_252_dout[29]),
  .I1(sdpb_inst_253_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3746 (
  .O(mux_o_3746),
  .I0(sdpb_inst_254_dout[29]),
  .I1(sdpb_inst_255_dout[29]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3747 (
  .O(mux_o_3747),
  .I0(mux_o_3683),
  .I1(mux_o_3684),
  .S0(dff_q_5)
);
MUX2 mux_inst_3748 (
  .O(mux_o_3748),
  .I0(mux_o_3685),
  .I1(mux_o_3686),
  .S0(dff_q_5)
);
MUX2 mux_inst_3749 (
  .O(mux_o_3749),
  .I0(mux_o_3687),
  .I1(mux_o_3688),
  .S0(dff_q_5)
);
MUX2 mux_inst_3750 (
  .O(mux_o_3750),
  .I0(mux_o_3689),
  .I1(mux_o_3690),
  .S0(dff_q_5)
);
MUX2 mux_inst_3751 (
  .O(mux_o_3751),
  .I0(mux_o_3691),
  .I1(mux_o_3692),
  .S0(dff_q_5)
);
MUX2 mux_inst_3752 (
  .O(mux_o_3752),
  .I0(mux_o_3693),
  .I1(mux_o_3694),
  .S0(dff_q_5)
);
MUX2 mux_inst_3753 (
  .O(mux_o_3753),
  .I0(mux_o_3695),
  .I1(mux_o_3696),
  .S0(dff_q_5)
);
MUX2 mux_inst_3754 (
  .O(mux_o_3754),
  .I0(mux_o_3697),
  .I1(mux_o_3698),
  .S0(dff_q_5)
);
MUX2 mux_inst_3755 (
  .O(mux_o_3755),
  .I0(mux_o_3699),
  .I1(mux_o_3700),
  .S0(dff_q_5)
);
MUX2 mux_inst_3756 (
  .O(mux_o_3756),
  .I0(mux_o_3701),
  .I1(mux_o_3702),
  .S0(dff_q_5)
);
MUX2 mux_inst_3757 (
  .O(mux_o_3757),
  .I0(mux_o_3703),
  .I1(mux_o_3704),
  .S0(dff_q_5)
);
MUX2 mux_inst_3758 (
  .O(mux_o_3758),
  .I0(mux_o_3705),
  .I1(mux_o_3706),
  .S0(dff_q_5)
);
MUX2 mux_inst_3759 (
  .O(mux_o_3759),
  .I0(mux_o_3707),
  .I1(mux_o_3708),
  .S0(dff_q_5)
);
MUX2 mux_inst_3760 (
  .O(mux_o_3760),
  .I0(mux_o_3709),
  .I1(mux_o_3710),
  .S0(dff_q_5)
);
MUX2 mux_inst_3761 (
  .O(mux_o_3761),
  .I0(mux_o_3711),
  .I1(mux_o_3712),
  .S0(dff_q_5)
);
MUX2 mux_inst_3762 (
  .O(mux_o_3762),
  .I0(mux_o_3713),
  .I1(mux_o_3714),
  .S0(dff_q_5)
);
MUX2 mux_inst_3763 (
  .O(mux_o_3763),
  .I0(mux_o_3715),
  .I1(mux_o_3716),
  .S0(dff_q_5)
);
MUX2 mux_inst_3764 (
  .O(mux_o_3764),
  .I0(mux_o_3717),
  .I1(mux_o_3718),
  .S0(dff_q_5)
);
MUX2 mux_inst_3765 (
  .O(mux_o_3765),
  .I0(mux_o_3719),
  .I1(mux_o_3720),
  .S0(dff_q_5)
);
MUX2 mux_inst_3766 (
  .O(mux_o_3766),
  .I0(mux_o_3721),
  .I1(mux_o_3722),
  .S0(dff_q_5)
);
MUX2 mux_inst_3767 (
  .O(mux_o_3767),
  .I0(mux_o_3723),
  .I1(mux_o_3724),
  .S0(dff_q_5)
);
MUX2 mux_inst_3768 (
  .O(mux_o_3768),
  .I0(mux_o_3725),
  .I1(mux_o_3726),
  .S0(dff_q_5)
);
MUX2 mux_inst_3769 (
  .O(mux_o_3769),
  .I0(mux_o_3727),
  .I1(mux_o_3728),
  .S0(dff_q_5)
);
MUX2 mux_inst_3770 (
  .O(mux_o_3770),
  .I0(mux_o_3729),
  .I1(mux_o_3730),
  .S0(dff_q_5)
);
MUX2 mux_inst_3771 (
  .O(mux_o_3771),
  .I0(mux_o_3731),
  .I1(mux_o_3732),
  .S0(dff_q_5)
);
MUX2 mux_inst_3772 (
  .O(mux_o_3772),
  .I0(mux_o_3733),
  .I1(mux_o_3734),
  .S0(dff_q_5)
);
MUX2 mux_inst_3773 (
  .O(mux_o_3773),
  .I0(mux_o_3735),
  .I1(mux_o_3736),
  .S0(dff_q_5)
);
MUX2 mux_inst_3774 (
  .O(mux_o_3774),
  .I0(mux_o_3737),
  .I1(mux_o_3738),
  .S0(dff_q_5)
);
MUX2 mux_inst_3775 (
  .O(mux_o_3775),
  .I0(mux_o_3739),
  .I1(mux_o_3740),
  .S0(dff_q_5)
);
MUX2 mux_inst_3776 (
  .O(mux_o_3776),
  .I0(mux_o_3741),
  .I1(mux_o_3742),
  .S0(dff_q_5)
);
MUX2 mux_inst_3777 (
  .O(mux_o_3777),
  .I0(mux_o_3743),
  .I1(mux_o_3744),
  .S0(dff_q_5)
);
MUX2 mux_inst_3778 (
  .O(mux_o_3778),
  .I0(mux_o_3745),
  .I1(mux_o_3746),
  .S0(dff_q_5)
);
MUX2 mux_inst_3779 (
  .O(mux_o_3779),
  .I0(mux_o_3747),
  .I1(mux_o_3748),
  .S0(dff_q_4)
);
MUX2 mux_inst_3780 (
  .O(mux_o_3780),
  .I0(mux_o_3749),
  .I1(mux_o_3750),
  .S0(dff_q_4)
);
MUX2 mux_inst_3781 (
  .O(mux_o_3781),
  .I0(mux_o_3751),
  .I1(mux_o_3752),
  .S0(dff_q_4)
);
MUX2 mux_inst_3782 (
  .O(mux_o_3782),
  .I0(mux_o_3753),
  .I1(mux_o_3754),
  .S0(dff_q_4)
);
MUX2 mux_inst_3783 (
  .O(mux_o_3783),
  .I0(mux_o_3755),
  .I1(mux_o_3756),
  .S0(dff_q_4)
);
MUX2 mux_inst_3784 (
  .O(mux_o_3784),
  .I0(mux_o_3757),
  .I1(mux_o_3758),
  .S0(dff_q_4)
);
MUX2 mux_inst_3785 (
  .O(mux_o_3785),
  .I0(mux_o_3759),
  .I1(mux_o_3760),
  .S0(dff_q_4)
);
MUX2 mux_inst_3786 (
  .O(mux_o_3786),
  .I0(mux_o_3761),
  .I1(mux_o_3762),
  .S0(dff_q_4)
);
MUX2 mux_inst_3787 (
  .O(mux_o_3787),
  .I0(mux_o_3763),
  .I1(mux_o_3764),
  .S0(dff_q_4)
);
MUX2 mux_inst_3788 (
  .O(mux_o_3788),
  .I0(mux_o_3765),
  .I1(mux_o_3766),
  .S0(dff_q_4)
);
MUX2 mux_inst_3789 (
  .O(mux_o_3789),
  .I0(mux_o_3767),
  .I1(mux_o_3768),
  .S0(dff_q_4)
);
MUX2 mux_inst_3790 (
  .O(mux_o_3790),
  .I0(mux_o_3769),
  .I1(mux_o_3770),
  .S0(dff_q_4)
);
MUX2 mux_inst_3791 (
  .O(mux_o_3791),
  .I0(mux_o_3771),
  .I1(mux_o_3772),
  .S0(dff_q_4)
);
MUX2 mux_inst_3792 (
  .O(mux_o_3792),
  .I0(mux_o_3773),
  .I1(mux_o_3774),
  .S0(dff_q_4)
);
MUX2 mux_inst_3793 (
  .O(mux_o_3793),
  .I0(mux_o_3775),
  .I1(mux_o_3776),
  .S0(dff_q_4)
);
MUX2 mux_inst_3794 (
  .O(mux_o_3794),
  .I0(mux_o_3777),
  .I1(mux_o_3778),
  .S0(dff_q_4)
);
MUX2 mux_inst_3795 (
  .O(mux_o_3795),
  .I0(mux_o_3779),
  .I1(mux_o_3780),
  .S0(dff_q_3)
);
MUX2 mux_inst_3796 (
  .O(mux_o_3796),
  .I0(mux_o_3781),
  .I1(mux_o_3782),
  .S0(dff_q_3)
);
MUX2 mux_inst_3797 (
  .O(mux_o_3797),
  .I0(mux_o_3783),
  .I1(mux_o_3784),
  .S0(dff_q_3)
);
MUX2 mux_inst_3798 (
  .O(mux_o_3798),
  .I0(mux_o_3785),
  .I1(mux_o_3786),
  .S0(dff_q_3)
);
MUX2 mux_inst_3799 (
  .O(mux_o_3799),
  .I0(mux_o_3787),
  .I1(mux_o_3788),
  .S0(dff_q_3)
);
MUX2 mux_inst_3800 (
  .O(mux_o_3800),
  .I0(mux_o_3789),
  .I1(mux_o_3790),
  .S0(dff_q_3)
);
MUX2 mux_inst_3801 (
  .O(mux_o_3801),
  .I0(mux_o_3791),
  .I1(mux_o_3792),
  .S0(dff_q_3)
);
MUX2 mux_inst_3802 (
  .O(mux_o_3802),
  .I0(mux_o_3793),
  .I1(mux_o_3794),
  .S0(dff_q_3)
);
MUX2 mux_inst_3803 (
  .O(mux_o_3803),
  .I0(mux_o_3795),
  .I1(mux_o_3796),
  .S0(dff_q_2)
);
MUX2 mux_inst_3804 (
  .O(mux_o_3804),
  .I0(mux_o_3797),
  .I1(mux_o_3798),
  .S0(dff_q_2)
);
MUX2 mux_inst_3805 (
  .O(mux_o_3805),
  .I0(mux_o_3799),
  .I1(mux_o_3800),
  .S0(dff_q_2)
);
MUX2 mux_inst_3806 (
  .O(mux_o_3806),
  .I0(mux_o_3801),
  .I1(mux_o_3802),
  .S0(dff_q_2)
);
MUX2 mux_inst_3807 (
  .O(mux_o_3807),
  .I0(mux_o_3803),
  .I1(mux_o_3804),
  .S0(dff_q_1)
);
MUX2 mux_inst_3808 (
  .O(mux_o_3808),
  .I0(mux_o_3805),
  .I1(mux_o_3806),
  .S0(dff_q_1)
);
MUX2 mux_inst_3809 (
  .O(dout[29]),
  .I0(mux_o_3807),
  .I1(mux_o_3808),
  .S0(dff_q_0)
);
MUX2 mux_inst_3810 (
  .O(mux_o_3810),
  .I0(sdpb_inst_128_dout[30]),
  .I1(sdpb_inst_129_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3811 (
  .O(mux_o_3811),
  .I0(sdpb_inst_130_dout[30]),
  .I1(sdpb_inst_131_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3812 (
  .O(mux_o_3812),
  .I0(sdpb_inst_132_dout[30]),
  .I1(sdpb_inst_133_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3813 (
  .O(mux_o_3813),
  .I0(sdpb_inst_134_dout[30]),
  .I1(sdpb_inst_135_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3814 (
  .O(mux_o_3814),
  .I0(sdpb_inst_136_dout[30]),
  .I1(sdpb_inst_137_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3815 (
  .O(mux_o_3815),
  .I0(sdpb_inst_138_dout[30]),
  .I1(sdpb_inst_139_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3816 (
  .O(mux_o_3816),
  .I0(sdpb_inst_140_dout[30]),
  .I1(sdpb_inst_141_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3817 (
  .O(mux_o_3817),
  .I0(sdpb_inst_142_dout[30]),
  .I1(sdpb_inst_143_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3818 (
  .O(mux_o_3818),
  .I0(sdpb_inst_144_dout[30]),
  .I1(sdpb_inst_145_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3819 (
  .O(mux_o_3819),
  .I0(sdpb_inst_146_dout[30]),
  .I1(sdpb_inst_147_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3820 (
  .O(mux_o_3820),
  .I0(sdpb_inst_148_dout[30]),
  .I1(sdpb_inst_149_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3821 (
  .O(mux_o_3821),
  .I0(sdpb_inst_150_dout[30]),
  .I1(sdpb_inst_151_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3822 (
  .O(mux_o_3822),
  .I0(sdpb_inst_152_dout[30]),
  .I1(sdpb_inst_153_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3823 (
  .O(mux_o_3823),
  .I0(sdpb_inst_154_dout[30]),
  .I1(sdpb_inst_155_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3824 (
  .O(mux_o_3824),
  .I0(sdpb_inst_156_dout[30]),
  .I1(sdpb_inst_157_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3825 (
  .O(mux_o_3825),
  .I0(sdpb_inst_158_dout[30]),
  .I1(sdpb_inst_159_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3826 (
  .O(mux_o_3826),
  .I0(sdpb_inst_160_dout[30]),
  .I1(sdpb_inst_161_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3827 (
  .O(mux_o_3827),
  .I0(sdpb_inst_162_dout[30]),
  .I1(sdpb_inst_163_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3828 (
  .O(mux_o_3828),
  .I0(sdpb_inst_164_dout[30]),
  .I1(sdpb_inst_165_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3829 (
  .O(mux_o_3829),
  .I0(sdpb_inst_166_dout[30]),
  .I1(sdpb_inst_167_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3830 (
  .O(mux_o_3830),
  .I0(sdpb_inst_168_dout[30]),
  .I1(sdpb_inst_169_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3831 (
  .O(mux_o_3831),
  .I0(sdpb_inst_170_dout[30]),
  .I1(sdpb_inst_171_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3832 (
  .O(mux_o_3832),
  .I0(sdpb_inst_172_dout[30]),
  .I1(sdpb_inst_173_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3833 (
  .O(mux_o_3833),
  .I0(sdpb_inst_174_dout[30]),
  .I1(sdpb_inst_175_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3834 (
  .O(mux_o_3834),
  .I0(sdpb_inst_176_dout[30]),
  .I1(sdpb_inst_177_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3835 (
  .O(mux_o_3835),
  .I0(sdpb_inst_178_dout[30]),
  .I1(sdpb_inst_179_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3836 (
  .O(mux_o_3836),
  .I0(sdpb_inst_180_dout[30]),
  .I1(sdpb_inst_181_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3837 (
  .O(mux_o_3837),
  .I0(sdpb_inst_182_dout[30]),
  .I1(sdpb_inst_183_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3838 (
  .O(mux_o_3838),
  .I0(sdpb_inst_184_dout[30]),
  .I1(sdpb_inst_185_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3839 (
  .O(mux_o_3839),
  .I0(sdpb_inst_186_dout[30]),
  .I1(sdpb_inst_187_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3840 (
  .O(mux_o_3840),
  .I0(sdpb_inst_188_dout[30]),
  .I1(sdpb_inst_189_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3841 (
  .O(mux_o_3841),
  .I0(sdpb_inst_190_dout[30]),
  .I1(sdpb_inst_191_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3842 (
  .O(mux_o_3842),
  .I0(sdpb_inst_192_dout[30]),
  .I1(sdpb_inst_193_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3843 (
  .O(mux_o_3843),
  .I0(sdpb_inst_194_dout[30]),
  .I1(sdpb_inst_195_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3844 (
  .O(mux_o_3844),
  .I0(sdpb_inst_196_dout[30]),
  .I1(sdpb_inst_197_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3845 (
  .O(mux_o_3845),
  .I0(sdpb_inst_198_dout[30]),
  .I1(sdpb_inst_199_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3846 (
  .O(mux_o_3846),
  .I0(sdpb_inst_200_dout[30]),
  .I1(sdpb_inst_201_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3847 (
  .O(mux_o_3847),
  .I0(sdpb_inst_202_dout[30]),
  .I1(sdpb_inst_203_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3848 (
  .O(mux_o_3848),
  .I0(sdpb_inst_204_dout[30]),
  .I1(sdpb_inst_205_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3849 (
  .O(mux_o_3849),
  .I0(sdpb_inst_206_dout[30]),
  .I1(sdpb_inst_207_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3850 (
  .O(mux_o_3850),
  .I0(sdpb_inst_208_dout[30]),
  .I1(sdpb_inst_209_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3851 (
  .O(mux_o_3851),
  .I0(sdpb_inst_210_dout[30]),
  .I1(sdpb_inst_211_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3852 (
  .O(mux_o_3852),
  .I0(sdpb_inst_212_dout[30]),
  .I1(sdpb_inst_213_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3853 (
  .O(mux_o_3853),
  .I0(sdpb_inst_214_dout[30]),
  .I1(sdpb_inst_215_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3854 (
  .O(mux_o_3854),
  .I0(sdpb_inst_216_dout[30]),
  .I1(sdpb_inst_217_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3855 (
  .O(mux_o_3855),
  .I0(sdpb_inst_218_dout[30]),
  .I1(sdpb_inst_219_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3856 (
  .O(mux_o_3856),
  .I0(sdpb_inst_220_dout[30]),
  .I1(sdpb_inst_221_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3857 (
  .O(mux_o_3857),
  .I0(sdpb_inst_222_dout[30]),
  .I1(sdpb_inst_223_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3858 (
  .O(mux_o_3858),
  .I0(sdpb_inst_224_dout[30]),
  .I1(sdpb_inst_225_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3859 (
  .O(mux_o_3859),
  .I0(sdpb_inst_226_dout[30]),
  .I1(sdpb_inst_227_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3860 (
  .O(mux_o_3860),
  .I0(sdpb_inst_228_dout[30]),
  .I1(sdpb_inst_229_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3861 (
  .O(mux_o_3861),
  .I0(sdpb_inst_230_dout[30]),
  .I1(sdpb_inst_231_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3862 (
  .O(mux_o_3862),
  .I0(sdpb_inst_232_dout[30]),
  .I1(sdpb_inst_233_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3863 (
  .O(mux_o_3863),
  .I0(sdpb_inst_234_dout[30]),
  .I1(sdpb_inst_235_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3864 (
  .O(mux_o_3864),
  .I0(sdpb_inst_236_dout[30]),
  .I1(sdpb_inst_237_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3865 (
  .O(mux_o_3865),
  .I0(sdpb_inst_238_dout[30]),
  .I1(sdpb_inst_239_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3866 (
  .O(mux_o_3866),
  .I0(sdpb_inst_240_dout[30]),
  .I1(sdpb_inst_241_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3867 (
  .O(mux_o_3867),
  .I0(sdpb_inst_242_dout[30]),
  .I1(sdpb_inst_243_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3868 (
  .O(mux_o_3868),
  .I0(sdpb_inst_244_dout[30]),
  .I1(sdpb_inst_245_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3869 (
  .O(mux_o_3869),
  .I0(sdpb_inst_246_dout[30]),
  .I1(sdpb_inst_247_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3870 (
  .O(mux_o_3870),
  .I0(sdpb_inst_248_dout[30]),
  .I1(sdpb_inst_249_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3871 (
  .O(mux_o_3871),
  .I0(sdpb_inst_250_dout[30]),
  .I1(sdpb_inst_251_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3872 (
  .O(mux_o_3872),
  .I0(sdpb_inst_252_dout[30]),
  .I1(sdpb_inst_253_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3873 (
  .O(mux_o_3873),
  .I0(sdpb_inst_254_dout[30]),
  .I1(sdpb_inst_255_dout[30]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3874 (
  .O(mux_o_3874),
  .I0(mux_o_3810),
  .I1(mux_o_3811),
  .S0(dff_q_5)
);
MUX2 mux_inst_3875 (
  .O(mux_o_3875),
  .I0(mux_o_3812),
  .I1(mux_o_3813),
  .S0(dff_q_5)
);
MUX2 mux_inst_3876 (
  .O(mux_o_3876),
  .I0(mux_o_3814),
  .I1(mux_o_3815),
  .S0(dff_q_5)
);
MUX2 mux_inst_3877 (
  .O(mux_o_3877),
  .I0(mux_o_3816),
  .I1(mux_o_3817),
  .S0(dff_q_5)
);
MUX2 mux_inst_3878 (
  .O(mux_o_3878),
  .I0(mux_o_3818),
  .I1(mux_o_3819),
  .S0(dff_q_5)
);
MUX2 mux_inst_3879 (
  .O(mux_o_3879),
  .I0(mux_o_3820),
  .I1(mux_o_3821),
  .S0(dff_q_5)
);
MUX2 mux_inst_3880 (
  .O(mux_o_3880),
  .I0(mux_o_3822),
  .I1(mux_o_3823),
  .S0(dff_q_5)
);
MUX2 mux_inst_3881 (
  .O(mux_o_3881),
  .I0(mux_o_3824),
  .I1(mux_o_3825),
  .S0(dff_q_5)
);
MUX2 mux_inst_3882 (
  .O(mux_o_3882),
  .I0(mux_o_3826),
  .I1(mux_o_3827),
  .S0(dff_q_5)
);
MUX2 mux_inst_3883 (
  .O(mux_o_3883),
  .I0(mux_o_3828),
  .I1(mux_o_3829),
  .S0(dff_q_5)
);
MUX2 mux_inst_3884 (
  .O(mux_o_3884),
  .I0(mux_o_3830),
  .I1(mux_o_3831),
  .S0(dff_q_5)
);
MUX2 mux_inst_3885 (
  .O(mux_o_3885),
  .I0(mux_o_3832),
  .I1(mux_o_3833),
  .S0(dff_q_5)
);
MUX2 mux_inst_3886 (
  .O(mux_o_3886),
  .I0(mux_o_3834),
  .I1(mux_o_3835),
  .S0(dff_q_5)
);
MUX2 mux_inst_3887 (
  .O(mux_o_3887),
  .I0(mux_o_3836),
  .I1(mux_o_3837),
  .S0(dff_q_5)
);
MUX2 mux_inst_3888 (
  .O(mux_o_3888),
  .I0(mux_o_3838),
  .I1(mux_o_3839),
  .S0(dff_q_5)
);
MUX2 mux_inst_3889 (
  .O(mux_o_3889),
  .I0(mux_o_3840),
  .I1(mux_o_3841),
  .S0(dff_q_5)
);
MUX2 mux_inst_3890 (
  .O(mux_o_3890),
  .I0(mux_o_3842),
  .I1(mux_o_3843),
  .S0(dff_q_5)
);
MUX2 mux_inst_3891 (
  .O(mux_o_3891),
  .I0(mux_o_3844),
  .I1(mux_o_3845),
  .S0(dff_q_5)
);
MUX2 mux_inst_3892 (
  .O(mux_o_3892),
  .I0(mux_o_3846),
  .I1(mux_o_3847),
  .S0(dff_q_5)
);
MUX2 mux_inst_3893 (
  .O(mux_o_3893),
  .I0(mux_o_3848),
  .I1(mux_o_3849),
  .S0(dff_q_5)
);
MUX2 mux_inst_3894 (
  .O(mux_o_3894),
  .I0(mux_o_3850),
  .I1(mux_o_3851),
  .S0(dff_q_5)
);
MUX2 mux_inst_3895 (
  .O(mux_o_3895),
  .I0(mux_o_3852),
  .I1(mux_o_3853),
  .S0(dff_q_5)
);
MUX2 mux_inst_3896 (
  .O(mux_o_3896),
  .I0(mux_o_3854),
  .I1(mux_o_3855),
  .S0(dff_q_5)
);
MUX2 mux_inst_3897 (
  .O(mux_o_3897),
  .I0(mux_o_3856),
  .I1(mux_o_3857),
  .S0(dff_q_5)
);
MUX2 mux_inst_3898 (
  .O(mux_o_3898),
  .I0(mux_o_3858),
  .I1(mux_o_3859),
  .S0(dff_q_5)
);
MUX2 mux_inst_3899 (
  .O(mux_o_3899),
  .I0(mux_o_3860),
  .I1(mux_o_3861),
  .S0(dff_q_5)
);
MUX2 mux_inst_3900 (
  .O(mux_o_3900),
  .I0(mux_o_3862),
  .I1(mux_o_3863),
  .S0(dff_q_5)
);
MUX2 mux_inst_3901 (
  .O(mux_o_3901),
  .I0(mux_o_3864),
  .I1(mux_o_3865),
  .S0(dff_q_5)
);
MUX2 mux_inst_3902 (
  .O(mux_o_3902),
  .I0(mux_o_3866),
  .I1(mux_o_3867),
  .S0(dff_q_5)
);
MUX2 mux_inst_3903 (
  .O(mux_o_3903),
  .I0(mux_o_3868),
  .I1(mux_o_3869),
  .S0(dff_q_5)
);
MUX2 mux_inst_3904 (
  .O(mux_o_3904),
  .I0(mux_o_3870),
  .I1(mux_o_3871),
  .S0(dff_q_5)
);
MUX2 mux_inst_3905 (
  .O(mux_o_3905),
  .I0(mux_o_3872),
  .I1(mux_o_3873),
  .S0(dff_q_5)
);
MUX2 mux_inst_3906 (
  .O(mux_o_3906),
  .I0(mux_o_3874),
  .I1(mux_o_3875),
  .S0(dff_q_4)
);
MUX2 mux_inst_3907 (
  .O(mux_o_3907),
  .I0(mux_o_3876),
  .I1(mux_o_3877),
  .S0(dff_q_4)
);
MUX2 mux_inst_3908 (
  .O(mux_o_3908),
  .I0(mux_o_3878),
  .I1(mux_o_3879),
  .S0(dff_q_4)
);
MUX2 mux_inst_3909 (
  .O(mux_o_3909),
  .I0(mux_o_3880),
  .I1(mux_o_3881),
  .S0(dff_q_4)
);
MUX2 mux_inst_3910 (
  .O(mux_o_3910),
  .I0(mux_o_3882),
  .I1(mux_o_3883),
  .S0(dff_q_4)
);
MUX2 mux_inst_3911 (
  .O(mux_o_3911),
  .I0(mux_o_3884),
  .I1(mux_o_3885),
  .S0(dff_q_4)
);
MUX2 mux_inst_3912 (
  .O(mux_o_3912),
  .I0(mux_o_3886),
  .I1(mux_o_3887),
  .S0(dff_q_4)
);
MUX2 mux_inst_3913 (
  .O(mux_o_3913),
  .I0(mux_o_3888),
  .I1(mux_o_3889),
  .S0(dff_q_4)
);
MUX2 mux_inst_3914 (
  .O(mux_o_3914),
  .I0(mux_o_3890),
  .I1(mux_o_3891),
  .S0(dff_q_4)
);
MUX2 mux_inst_3915 (
  .O(mux_o_3915),
  .I0(mux_o_3892),
  .I1(mux_o_3893),
  .S0(dff_q_4)
);
MUX2 mux_inst_3916 (
  .O(mux_o_3916),
  .I0(mux_o_3894),
  .I1(mux_o_3895),
  .S0(dff_q_4)
);
MUX2 mux_inst_3917 (
  .O(mux_o_3917),
  .I0(mux_o_3896),
  .I1(mux_o_3897),
  .S0(dff_q_4)
);
MUX2 mux_inst_3918 (
  .O(mux_o_3918),
  .I0(mux_o_3898),
  .I1(mux_o_3899),
  .S0(dff_q_4)
);
MUX2 mux_inst_3919 (
  .O(mux_o_3919),
  .I0(mux_o_3900),
  .I1(mux_o_3901),
  .S0(dff_q_4)
);
MUX2 mux_inst_3920 (
  .O(mux_o_3920),
  .I0(mux_o_3902),
  .I1(mux_o_3903),
  .S0(dff_q_4)
);
MUX2 mux_inst_3921 (
  .O(mux_o_3921),
  .I0(mux_o_3904),
  .I1(mux_o_3905),
  .S0(dff_q_4)
);
MUX2 mux_inst_3922 (
  .O(mux_o_3922),
  .I0(mux_o_3906),
  .I1(mux_o_3907),
  .S0(dff_q_3)
);
MUX2 mux_inst_3923 (
  .O(mux_o_3923),
  .I0(mux_o_3908),
  .I1(mux_o_3909),
  .S0(dff_q_3)
);
MUX2 mux_inst_3924 (
  .O(mux_o_3924),
  .I0(mux_o_3910),
  .I1(mux_o_3911),
  .S0(dff_q_3)
);
MUX2 mux_inst_3925 (
  .O(mux_o_3925),
  .I0(mux_o_3912),
  .I1(mux_o_3913),
  .S0(dff_q_3)
);
MUX2 mux_inst_3926 (
  .O(mux_o_3926),
  .I0(mux_o_3914),
  .I1(mux_o_3915),
  .S0(dff_q_3)
);
MUX2 mux_inst_3927 (
  .O(mux_o_3927),
  .I0(mux_o_3916),
  .I1(mux_o_3917),
  .S0(dff_q_3)
);
MUX2 mux_inst_3928 (
  .O(mux_o_3928),
  .I0(mux_o_3918),
  .I1(mux_o_3919),
  .S0(dff_q_3)
);
MUX2 mux_inst_3929 (
  .O(mux_o_3929),
  .I0(mux_o_3920),
  .I1(mux_o_3921),
  .S0(dff_q_3)
);
MUX2 mux_inst_3930 (
  .O(mux_o_3930),
  .I0(mux_o_3922),
  .I1(mux_o_3923),
  .S0(dff_q_2)
);
MUX2 mux_inst_3931 (
  .O(mux_o_3931),
  .I0(mux_o_3924),
  .I1(mux_o_3925),
  .S0(dff_q_2)
);
MUX2 mux_inst_3932 (
  .O(mux_o_3932),
  .I0(mux_o_3926),
  .I1(mux_o_3927),
  .S0(dff_q_2)
);
MUX2 mux_inst_3933 (
  .O(mux_o_3933),
  .I0(mux_o_3928),
  .I1(mux_o_3929),
  .S0(dff_q_2)
);
MUX2 mux_inst_3934 (
  .O(mux_o_3934),
  .I0(mux_o_3930),
  .I1(mux_o_3931),
  .S0(dff_q_1)
);
MUX2 mux_inst_3935 (
  .O(mux_o_3935),
  .I0(mux_o_3932),
  .I1(mux_o_3933),
  .S0(dff_q_1)
);
MUX2 mux_inst_3936 (
  .O(dout[30]),
  .I0(mux_o_3934),
  .I1(mux_o_3935),
  .S0(dff_q_0)
);
MUX2 mux_inst_3937 (
  .O(mux_o_3937),
  .I0(sdpb_inst_128_dout[31]),
  .I1(sdpb_inst_129_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3938 (
  .O(mux_o_3938),
  .I0(sdpb_inst_130_dout[31]),
  .I1(sdpb_inst_131_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3939 (
  .O(mux_o_3939),
  .I0(sdpb_inst_132_dout[31]),
  .I1(sdpb_inst_133_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3940 (
  .O(mux_o_3940),
  .I0(sdpb_inst_134_dout[31]),
  .I1(sdpb_inst_135_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3941 (
  .O(mux_o_3941),
  .I0(sdpb_inst_136_dout[31]),
  .I1(sdpb_inst_137_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3942 (
  .O(mux_o_3942),
  .I0(sdpb_inst_138_dout[31]),
  .I1(sdpb_inst_139_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3943 (
  .O(mux_o_3943),
  .I0(sdpb_inst_140_dout[31]),
  .I1(sdpb_inst_141_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3944 (
  .O(mux_o_3944),
  .I0(sdpb_inst_142_dout[31]),
  .I1(sdpb_inst_143_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3945 (
  .O(mux_o_3945),
  .I0(sdpb_inst_144_dout[31]),
  .I1(sdpb_inst_145_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3946 (
  .O(mux_o_3946),
  .I0(sdpb_inst_146_dout[31]),
  .I1(sdpb_inst_147_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3947 (
  .O(mux_o_3947),
  .I0(sdpb_inst_148_dout[31]),
  .I1(sdpb_inst_149_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3948 (
  .O(mux_o_3948),
  .I0(sdpb_inst_150_dout[31]),
  .I1(sdpb_inst_151_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3949 (
  .O(mux_o_3949),
  .I0(sdpb_inst_152_dout[31]),
  .I1(sdpb_inst_153_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3950 (
  .O(mux_o_3950),
  .I0(sdpb_inst_154_dout[31]),
  .I1(sdpb_inst_155_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3951 (
  .O(mux_o_3951),
  .I0(sdpb_inst_156_dout[31]),
  .I1(sdpb_inst_157_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3952 (
  .O(mux_o_3952),
  .I0(sdpb_inst_158_dout[31]),
  .I1(sdpb_inst_159_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3953 (
  .O(mux_o_3953),
  .I0(sdpb_inst_160_dout[31]),
  .I1(sdpb_inst_161_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3954 (
  .O(mux_o_3954),
  .I0(sdpb_inst_162_dout[31]),
  .I1(sdpb_inst_163_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3955 (
  .O(mux_o_3955),
  .I0(sdpb_inst_164_dout[31]),
  .I1(sdpb_inst_165_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3956 (
  .O(mux_o_3956),
  .I0(sdpb_inst_166_dout[31]),
  .I1(sdpb_inst_167_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3957 (
  .O(mux_o_3957),
  .I0(sdpb_inst_168_dout[31]),
  .I1(sdpb_inst_169_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3958 (
  .O(mux_o_3958),
  .I0(sdpb_inst_170_dout[31]),
  .I1(sdpb_inst_171_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3959 (
  .O(mux_o_3959),
  .I0(sdpb_inst_172_dout[31]),
  .I1(sdpb_inst_173_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3960 (
  .O(mux_o_3960),
  .I0(sdpb_inst_174_dout[31]),
  .I1(sdpb_inst_175_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3961 (
  .O(mux_o_3961),
  .I0(sdpb_inst_176_dout[31]),
  .I1(sdpb_inst_177_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3962 (
  .O(mux_o_3962),
  .I0(sdpb_inst_178_dout[31]),
  .I1(sdpb_inst_179_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3963 (
  .O(mux_o_3963),
  .I0(sdpb_inst_180_dout[31]),
  .I1(sdpb_inst_181_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3964 (
  .O(mux_o_3964),
  .I0(sdpb_inst_182_dout[31]),
  .I1(sdpb_inst_183_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3965 (
  .O(mux_o_3965),
  .I0(sdpb_inst_184_dout[31]),
  .I1(sdpb_inst_185_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3966 (
  .O(mux_o_3966),
  .I0(sdpb_inst_186_dout[31]),
  .I1(sdpb_inst_187_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3967 (
  .O(mux_o_3967),
  .I0(sdpb_inst_188_dout[31]),
  .I1(sdpb_inst_189_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3968 (
  .O(mux_o_3968),
  .I0(sdpb_inst_190_dout[31]),
  .I1(sdpb_inst_191_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3969 (
  .O(mux_o_3969),
  .I0(sdpb_inst_192_dout[31]),
  .I1(sdpb_inst_193_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3970 (
  .O(mux_o_3970),
  .I0(sdpb_inst_194_dout[31]),
  .I1(sdpb_inst_195_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3971 (
  .O(mux_o_3971),
  .I0(sdpb_inst_196_dout[31]),
  .I1(sdpb_inst_197_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3972 (
  .O(mux_o_3972),
  .I0(sdpb_inst_198_dout[31]),
  .I1(sdpb_inst_199_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3973 (
  .O(mux_o_3973),
  .I0(sdpb_inst_200_dout[31]),
  .I1(sdpb_inst_201_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3974 (
  .O(mux_o_3974),
  .I0(sdpb_inst_202_dout[31]),
  .I1(sdpb_inst_203_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3975 (
  .O(mux_o_3975),
  .I0(sdpb_inst_204_dout[31]),
  .I1(sdpb_inst_205_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3976 (
  .O(mux_o_3976),
  .I0(sdpb_inst_206_dout[31]),
  .I1(sdpb_inst_207_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3977 (
  .O(mux_o_3977),
  .I0(sdpb_inst_208_dout[31]),
  .I1(sdpb_inst_209_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3978 (
  .O(mux_o_3978),
  .I0(sdpb_inst_210_dout[31]),
  .I1(sdpb_inst_211_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3979 (
  .O(mux_o_3979),
  .I0(sdpb_inst_212_dout[31]),
  .I1(sdpb_inst_213_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3980 (
  .O(mux_o_3980),
  .I0(sdpb_inst_214_dout[31]),
  .I1(sdpb_inst_215_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3981 (
  .O(mux_o_3981),
  .I0(sdpb_inst_216_dout[31]),
  .I1(sdpb_inst_217_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3982 (
  .O(mux_o_3982),
  .I0(sdpb_inst_218_dout[31]),
  .I1(sdpb_inst_219_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3983 (
  .O(mux_o_3983),
  .I0(sdpb_inst_220_dout[31]),
  .I1(sdpb_inst_221_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3984 (
  .O(mux_o_3984),
  .I0(sdpb_inst_222_dout[31]),
  .I1(sdpb_inst_223_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3985 (
  .O(mux_o_3985),
  .I0(sdpb_inst_224_dout[31]),
  .I1(sdpb_inst_225_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3986 (
  .O(mux_o_3986),
  .I0(sdpb_inst_226_dout[31]),
  .I1(sdpb_inst_227_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3987 (
  .O(mux_o_3987),
  .I0(sdpb_inst_228_dout[31]),
  .I1(sdpb_inst_229_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3988 (
  .O(mux_o_3988),
  .I0(sdpb_inst_230_dout[31]),
  .I1(sdpb_inst_231_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3989 (
  .O(mux_o_3989),
  .I0(sdpb_inst_232_dout[31]),
  .I1(sdpb_inst_233_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3990 (
  .O(mux_o_3990),
  .I0(sdpb_inst_234_dout[31]),
  .I1(sdpb_inst_235_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3991 (
  .O(mux_o_3991),
  .I0(sdpb_inst_236_dout[31]),
  .I1(sdpb_inst_237_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3992 (
  .O(mux_o_3992),
  .I0(sdpb_inst_238_dout[31]),
  .I1(sdpb_inst_239_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3993 (
  .O(mux_o_3993),
  .I0(sdpb_inst_240_dout[31]),
  .I1(sdpb_inst_241_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3994 (
  .O(mux_o_3994),
  .I0(sdpb_inst_242_dout[31]),
  .I1(sdpb_inst_243_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3995 (
  .O(mux_o_3995),
  .I0(sdpb_inst_244_dout[31]),
  .I1(sdpb_inst_245_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3996 (
  .O(mux_o_3996),
  .I0(sdpb_inst_246_dout[31]),
  .I1(sdpb_inst_247_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3997 (
  .O(mux_o_3997),
  .I0(sdpb_inst_248_dout[31]),
  .I1(sdpb_inst_249_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3998 (
  .O(mux_o_3998),
  .I0(sdpb_inst_250_dout[31]),
  .I1(sdpb_inst_251_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_3999 (
  .O(mux_o_3999),
  .I0(sdpb_inst_252_dout[31]),
  .I1(sdpb_inst_253_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_4000 (
  .O(mux_o_4000),
  .I0(sdpb_inst_254_dout[31]),
  .I1(sdpb_inst_255_dout[31]),
  .S0(dff_q_6)
);
MUX2 mux_inst_4001 (
  .O(mux_o_4001),
  .I0(mux_o_3937),
  .I1(mux_o_3938),
  .S0(dff_q_5)
);
MUX2 mux_inst_4002 (
  .O(mux_o_4002),
  .I0(mux_o_3939),
  .I1(mux_o_3940),
  .S0(dff_q_5)
);
MUX2 mux_inst_4003 (
  .O(mux_o_4003),
  .I0(mux_o_3941),
  .I1(mux_o_3942),
  .S0(dff_q_5)
);
MUX2 mux_inst_4004 (
  .O(mux_o_4004),
  .I0(mux_o_3943),
  .I1(mux_o_3944),
  .S0(dff_q_5)
);
MUX2 mux_inst_4005 (
  .O(mux_o_4005),
  .I0(mux_o_3945),
  .I1(mux_o_3946),
  .S0(dff_q_5)
);
MUX2 mux_inst_4006 (
  .O(mux_o_4006),
  .I0(mux_o_3947),
  .I1(mux_o_3948),
  .S0(dff_q_5)
);
MUX2 mux_inst_4007 (
  .O(mux_o_4007),
  .I0(mux_o_3949),
  .I1(mux_o_3950),
  .S0(dff_q_5)
);
MUX2 mux_inst_4008 (
  .O(mux_o_4008),
  .I0(mux_o_3951),
  .I1(mux_o_3952),
  .S0(dff_q_5)
);
MUX2 mux_inst_4009 (
  .O(mux_o_4009),
  .I0(mux_o_3953),
  .I1(mux_o_3954),
  .S0(dff_q_5)
);
MUX2 mux_inst_4010 (
  .O(mux_o_4010),
  .I0(mux_o_3955),
  .I1(mux_o_3956),
  .S0(dff_q_5)
);
MUX2 mux_inst_4011 (
  .O(mux_o_4011),
  .I0(mux_o_3957),
  .I1(mux_o_3958),
  .S0(dff_q_5)
);
MUX2 mux_inst_4012 (
  .O(mux_o_4012),
  .I0(mux_o_3959),
  .I1(mux_o_3960),
  .S0(dff_q_5)
);
MUX2 mux_inst_4013 (
  .O(mux_o_4013),
  .I0(mux_o_3961),
  .I1(mux_o_3962),
  .S0(dff_q_5)
);
MUX2 mux_inst_4014 (
  .O(mux_o_4014),
  .I0(mux_o_3963),
  .I1(mux_o_3964),
  .S0(dff_q_5)
);
MUX2 mux_inst_4015 (
  .O(mux_o_4015),
  .I0(mux_o_3965),
  .I1(mux_o_3966),
  .S0(dff_q_5)
);
MUX2 mux_inst_4016 (
  .O(mux_o_4016),
  .I0(mux_o_3967),
  .I1(mux_o_3968),
  .S0(dff_q_5)
);
MUX2 mux_inst_4017 (
  .O(mux_o_4017),
  .I0(mux_o_3969),
  .I1(mux_o_3970),
  .S0(dff_q_5)
);
MUX2 mux_inst_4018 (
  .O(mux_o_4018),
  .I0(mux_o_3971),
  .I1(mux_o_3972),
  .S0(dff_q_5)
);
MUX2 mux_inst_4019 (
  .O(mux_o_4019),
  .I0(mux_o_3973),
  .I1(mux_o_3974),
  .S0(dff_q_5)
);
MUX2 mux_inst_4020 (
  .O(mux_o_4020),
  .I0(mux_o_3975),
  .I1(mux_o_3976),
  .S0(dff_q_5)
);
MUX2 mux_inst_4021 (
  .O(mux_o_4021),
  .I0(mux_o_3977),
  .I1(mux_o_3978),
  .S0(dff_q_5)
);
MUX2 mux_inst_4022 (
  .O(mux_o_4022),
  .I0(mux_o_3979),
  .I1(mux_o_3980),
  .S0(dff_q_5)
);
MUX2 mux_inst_4023 (
  .O(mux_o_4023),
  .I0(mux_o_3981),
  .I1(mux_o_3982),
  .S0(dff_q_5)
);
MUX2 mux_inst_4024 (
  .O(mux_o_4024),
  .I0(mux_o_3983),
  .I1(mux_o_3984),
  .S0(dff_q_5)
);
MUX2 mux_inst_4025 (
  .O(mux_o_4025),
  .I0(mux_o_3985),
  .I1(mux_o_3986),
  .S0(dff_q_5)
);
MUX2 mux_inst_4026 (
  .O(mux_o_4026),
  .I0(mux_o_3987),
  .I1(mux_o_3988),
  .S0(dff_q_5)
);
MUX2 mux_inst_4027 (
  .O(mux_o_4027),
  .I0(mux_o_3989),
  .I1(mux_o_3990),
  .S0(dff_q_5)
);
MUX2 mux_inst_4028 (
  .O(mux_o_4028),
  .I0(mux_o_3991),
  .I1(mux_o_3992),
  .S0(dff_q_5)
);
MUX2 mux_inst_4029 (
  .O(mux_o_4029),
  .I0(mux_o_3993),
  .I1(mux_o_3994),
  .S0(dff_q_5)
);
MUX2 mux_inst_4030 (
  .O(mux_o_4030),
  .I0(mux_o_3995),
  .I1(mux_o_3996),
  .S0(dff_q_5)
);
MUX2 mux_inst_4031 (
  .O(mux_o_4031),
  .I0(mux_o_3997),
  .I1(mux_o_3998),
  .S0(dff_q_5)
);
MUX2 mux_inst_4032 (
  .O(mux_o_4032),
  .I0(mux_o_3999),
  .I1(mux_o_4000),
  .S0(dff_q_5)
);
MUX2 mux_inst_4033 (
  .O(mux_o_4033),
  .I0(mux_o_4001),
  .I1(mux_o_4002),
  .S0(dff_q_4)
);
MUX2 mux_inst_4034 (
  .O(mux_o_4034),
  .I0(mux_o_4003),
  .I1(mux_o_4004),
  .S0(dff_q_4)
);
MUX2 mux_inst_4035 (
  .O(mux_o_4035),
  .I0(mux_o_4005),
  .I1(mux_o_4006),
  .S0(dff_q_4)
);
MUX2 mux_inst_4036 (
  .O(mux_o_4036),
  .I0(mux_o_4007),
  .I1(mux_o_4008),
  .S0(dff_q_4)
);
MUX2 mux_inst_4037 (
  .O(mux_o_4037),
  .I0(mux_o_4009),
  .I1(mux_o_4010),
  .S0(dff_q_4)
);
MUX2 mux_inst_4038 (
  .O(mux_o_4038),
  .I0(mux_o_4011),
  .I1(mux_o_4012),
  .S0(dff_q_4)
);
MUX2 mux_inst_4039 (
  .O(mux_o_4039),
  .I0(mux_o_4013),
  .I1(mux_o_4014),
  .S0(dff_q_4)
);
MUX2 mux_inst_4040 (
  .O(mux_o_4040),
  .I0(mux_o_4015),
  .I1(mux_o_4016),
  .S0(dff_q_4)
);
MUX2 mux_inst_4041 (
  .O(mux_o_4041),
  .I0(mux_o_4017),
  .I1(mux_o_4018),
  .S0(dff_q_4)
);
MUX2 mux_inst_4042 (
  .O(mux_o_4042),
  .I0(mux_o_4019),
  .I1(mux_o_4020),
  .S0(dff_q_4)
);
MUX2 mux_inst_4043 (
  .O(mux_o_4043),
  .I0(mux_o_4021),
  .I1(mux_o_4022),
  .S0(dff_q_4)
);
MUX2 mux_inst_4044 (
  .O(mux_o_4044),
  .I0(mux_o_4023),
  .I1(mux_o_4024),
  .S0(dff_q_4)
);
MUX2 mux_inst_4045 (
  .O(mux_o_4045),
  .I0(mux_o_4025),
  .I1(mux_o_4026),
  .S0(dff_q_4)
);
MUX2 mux_inst_4046 (
  .O(mux_o_4046),
  .I0(mux_o_4027),
  .I1(mux_o_4028),
  .S0(dff_q_4)
);
MUX2 mux_inst_4047 (
  .O(mux_o_4047),
  .I0(mux_o_4029),
  .I1(mux_o_4030),
  .S0(dff_q_4)
);
MUX2 mux_inst_4048 (
  .O(mux_o_4048),
  .I0(mux_o_4031),
  .I1(mux_o_4032),
  .S0(dff_q_4)
);
MUX2 mux_inst_4049 (
  .O(mux_o_4049),
  .I0(mux_o_4033),
  .I1(mux_o_4034),
  .S0(dff_q_3)
);
MUX2 mux_inst_4050 (
  .O(mux_o_4050),
  .I0(mux_o_4035),
  .I1(mux_o_4036),
  .S0(dff_q_3)
);
MUX2 mux_inst_4051 (
  .O(mux_o_4051),
  .I0(mux_o_4037),
  .I1(mux_o_4038),
  .S0(dff_q_3)
);
MUX2 mux_inst_4052 (
  .O(mux_o_4052),
  .I0(mux_o_4039),
  .I1(mux_o_4040),
  .S0(dff_q_3)
);
MUX2 mux_inst_4053 (
  .O(mux_o_4053),
  .I0(mux_o_4041),
  .I1(mux_o_4042),
  .S0(dff_q_3)
);
MUX2 mux_inst_4054 (
  .O(mux_o_4054),
  .I0(mux_o_4043),
  .I1(mux_o_4044),
  .S0(dff_q_3)
);
MUX2 mux_inst_4055 (
  .O(mux_o_4055),
  .I0(mux_o_4045),
  .I1(mux_o_4046),
  .S0(dff_q_3)
);
MUX2 mux_inst_4056 (
  .O(mux_o_4056),
  .I0(mux_o_4047),
  .I1(mux_o_4048),
  .S0(dff_q_3)
);
MUX2 mux_inst_4057 (
  .O(mux_o_4057),
  .I0(mux_o_4049),
  .I1(mux_o_4050),
  .S0(dff_q_2)
);
MUX2 mux_inst_4058 (
  .O(mux_o_4058),
  .I0(mux_o_4051),
  .I1(mux_o_4052),
  .S0(dff_q_2)
);
MUX2 mux_inst_4059 (
  .O(mux_o_4059),
  .I0(mux_o_4053),
  .I1(mux_o_4054),
  .S0(dff_q_2)
);
MUX2 mux_inst_4060 (
  .O(mux_o_4060),
  .I0(mux_o_4055),
  .I1(mux_o_4056),
  .S0(dff_q_2)
);
MUX2 mux_inst_4061 (
  .O(mux_o_4061),
  .I0(mux_o_4057),
  .I1(mux_o_4058),
  .S0(dff_q_1)
);
MUX2 mux_inst_4062 (
  .O(mux_o_4062),
  .I0(mux_o_4059),
  .I1(mux_o_4060),
  .S0(dff_q_1)
);
MUX2 mux_inst_4063 (
  .O(dout[31]),
  .I0(mux_o_4061),
  .I1(mux_o_4062),
  .S0(dff_q_0)
);
endmodule //SRAM_SDPB
